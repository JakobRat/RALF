magic
tech sky130A
magscale 1 2
timestamp 1702632978
<< checkpaint >>
rect -1556 -1797 1556 1797
<< nwell >>
rect -296 -537 296 537
<< pmos >>
rect -100 118 100 318
rect -100 -318 100 -118
<< pdiff >>
rect -158 306 -100 318
rect -158 130 -146 306
rect -112 130 -100 306
rect -158 118 -100 130
rect 100 306 158 318
rect 100 130 112 306
rect 146 130 158 306
rect 100 118 158 130
rect -158 -130 -100 -118
rect -158 -306 -146 -130
rect -112 -306 -100 -130
rect -158 -318 -100 -306
rect 100 -130 158 -118
rect 100 -306 112 -130
rect 146 -306 158 -130
rect 100 -318 158 -306
<< pdiffc >>
rect -146 130 -112 306
rect 112 130 146 306
rect -146 -306 -112 -130
rect 112 -306 146 -130
<< nsubdiff >>
rect -260 467 260 501
rect -260 -467 -226 467
rect 226 -467 260 467
rect -260 -501 -164 -467
rect 164 -501 260 -467
<< nsubdiffcont >>
rect -164 -501 164 -467
<< poly >>
rect -100 399 100 415
rect -100 365 -84 399
rect 84 365 100 399
rect -100 318 100 365
rect -100 71 100 118
rect -100 37 -84 71
rect 84 37 100 71
rect -100 21 100 37
rect -100 -37 100 -21
rect -100 -71 -84 -37
rect 84 -71 100 -37
rect -100 -118 100 -71
rect -100 -365 100 -318
rect -100 -399 -84 -365
rect 84 -399 100 -365
rect -100 -415 100 -399
<< polycont >>
rect -84 365 84 399
rect -84 37 84 71
rect -84 -71 84 -37
rect -84 -399 84 -365
<< locali >>
rect -260 467 260 501
rect -260 -467 -226 467
rect -100 365 -84 399
rect 84 365 100 399
rect -146 306 -112 322
rect -146 114 -112 130
rect 112 306 146 322
rect 112 114 146 130
rect -100 37 -84 71
rect 84 37 100 71
rect -100 -71 -84 -37
rect 84 -71 100 -37
rect -146 -130 -112 -114
rect -146 -322 -112 -306
rect 112 -130 146 -114
rect 112 -322 146 -306
rect -100 -399 -84 -365
rect 84 -399 100 -365
rect 226 -467 260 467
rect -260 -501 -164 -467
rect 164 -501 260 -467
<< properties >>
string FIXED_BBOX -243 -484 243 484
<< end >>
