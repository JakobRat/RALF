** sch_path: /home/jakob/Documents/AutomatedLayoutGeneration/Circuits/MillerOpAmp/MillerOpAmp.sch
**.subckt MillerOpAmp Von Vop Vbias2 Vp Vn Vbias1 VPWR VGND
*.opin Von
*.opin Vop
*.ipin Vbias2
*.ipin Vp
*.ipin Vn
*.ipin Vbias1
*.iopin VPWR
*.iopin VGND
x1 VPWR Vbias2 Von1 Vop1 Vp Vn Vbias1 VGND DiffAmp
x2 VPWR Von1 Von Vbias1 VGND CSAmp
x3 VPWR Vop1 Vop Vbias1 VGND CSAmp
XC1 Von1 Von sky130_fd_pr__cap_mim_m3_1 W=5 L=5 MF=1 m=1
XC2 Vop1 Vop sky130_fd_pr__cap_mim_m3_1 W=5 L=5 MF=1 m=1
**.ends

* expanding   symbol:
*+  /home/jakob/Documents/AutomatedLayoutGeneration/Circuits/MillerOpAmp/DiffAmp.sym # of pins=8
** sym_path: /home/jakob/Documents/AutomatedLayoutGeneration/Circuits/MillerOpAmp/DiffAmp.sym
** sch_path: /home/jakob/Documents/AutomatedLayoutGeneration/Circuits/MillerOpAmp/DiffAmp.sch
.subckt DiffAmp Vdd Vbias2 Von Vop Vp Vn Vbias1 Vss
*.iopin Vdd
*.iopin Vss
*.ipin Vp
*.ipin Vn
*.ipin Vbias1
*.ipin Vbias2
*.opin Vop
*.opin Von
XM1 Vop Vp Vmid Vss sky130_fd_pr__nfet_01v8 L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM2 Von Vn Vmid Vss sky130_fd_pr__nfet_01v8 L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM3 Vop Vbias2 Vdd Vdd sky130_fd_pr__pfet_01v8 L=1 W=2 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM4 Von Vbias2 Vdd Vdd sky130_fd_pr__pfet_01v8 L=1 W=2 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM5 Vmid Vbias1 Vss Vss sky130_fd_pr__nfet_01v8 L=2 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:
*+  /home/jakob/Documents/AutomatedLayoutGeneration/Circuits/MillerOpAmp/CSAmp.sym # of pins=5
** sym_path: /home/jakob/Documents/AutomatedLayoutGeneration/Circuits/MillerOpAmp/CSAmp.sym
** sch_path: /home/jakob/Documents/AutomatedLayoutGeneration/Circuits/MillerOpAmp/CSAmp.sch
.subckt CSAmp Vdd Vi Vo Vbias1 Vss
*.ipin Vbias1
*.ipin Vi
*.iopin Vdd
*.iopin Vss
*.opin Vo
XM1 Vo Vi Vdd Vdd sky130_fd_pr__pfet_01v8 L=1 W=4 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM2 Vo Vbias1 Vss Vss sky130_fd_pr__nfet_01v8 L=2 W=8 nf=4 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
.ends

.end