magic
tech sky130A
magscale 1 2
timestamp 1701937426
<< checkpaint >>
rect -1876 -2033 1876 2033
<< pwell >>
rect -616 -773 616 773
<< psubdiff >>
rect -580 703 580 737
rect -580 -703 -546 703
rect 546 -703 580 703
rect -580 -737 -484 -703
rect 484 -737 580 -703
<< psubdiffcont >>
rect -484 -737 484 -703
<< xpolycontact >>
rect -450 175 -380 607
rect -450 -607 -380 -175
rect -284 175 -214 607
rect -284 -607 -214 -175
rect -118 175 -48 607
rect -118 -607 -48 -175
rect 48 175 118 607
rect 48 -607 118 -175
rect 214 175 284 607
rect 214 -607 284 -175
rect 380 175 450 607
rect 380 -607 450 -175
<< xpolyres >>
rect -450 -175 -380 175
rect -284 -175 -214 175
rect -118 -175 -48 175
rect 48 -175 118 175
rect 214 -175 284 175
rect 380 -175 450 175
<< locali >>
rect -500 -737 -484 -703
rect 484 -737 500 -703
<< res0p35 >>
rect -452 -177 -378 177
rect -286 -177 -212 177
rect -120 -177 -46 177
rect 46 -177 120 177
rect 212 -177 286 177
rect 378 -177 452 177
<< properties >>
string FIXED_BBOX -563 -720 563 720
<< end >>
