magic
tech sky130A
magscale 1 2
timestamp 1702720037
<< checkpaint >>
rect -303 2701 3067 2809
rect -1261 1797 3067 2701
rect -1556 1739 3067 1797
rect -1685 1685 3067 1739
rect -1739 1556 3067 1685
rect -1797 -669 3067 1556
rect -1797 -1261 2333 -669
rect -1797 -1556 1797 -1261
rect -1739 -1685 1739 -1556
rect -1685 -1739 1685 -1685
rect -1556 -1797 1556 -1739
use XCCP_XM3_XM4  XCCP_XM3_XM4_0 ~/Documents/RALF/Magic/Devices
timestamp 1702720036
transform 0 1 536 -1 0 295
box -296 -537 296 537
use XDP_XM1_XM2  XDP_XM1_XM2_0 ~/Documents/RALF/Magic/Devices
timestamp 1702720036
transform 0 -1 478 1 0 1016
box -425 -479 425 479
use XM5  XM5_0 ~/Documents/RALF/Magic/Devices
timestamp 1702720036
transform 1 0 1382 0 1 1070
box -425 -479 425 479
<< end >>
