magic
tech sky130A
magscale 1 2
timestamp 1702573428
<< checkpaint >>
rect -1656 -1539 1656 1539
<< pwell >>
rect -396 -279 396 279
<< nmos >>
rect -200 -131 200 69
<< ndiff >>
rect -258 57 -200 69
rect -258 -119 -246 57
rect -212 -119 -200 57
rect -258 -131 -200 -119
rect 200 57 258 69
rect 200 -119 212 57
rect 246 -119 258 57
rect 200 -131 258 -119
<< ndiffc >>
rect -246 -119 -212 57
rect 212 -119 246 57
<< psubdiff >>
rect -360 209 360 243
rect -360 -209 -326 209
rect 326 -209 360 209
rect -360 -243 -264 -209
rect 264 -243 360 -209
<< psubdiffcont >>
rect -264 -243 264 -209
<< poly >>
rect -200 141 200 157
rect -200 107 -184 141
rect 184 107 200 141
rect -200 69 200 107
rect -200 -157 200 -131
<< polycont >>
rect -184 107 184 141
<< locali >>
rect -360 209 360 243
rect -360 -209 -326 209
rect -200 107 -184 141
rect 184 107 200 141
rect -246 57 -212 73
rect -246 -135 -212 -119
rect 212 57 246 73
rect 212 -135 246 -119
rect 326 -209 360 209
rect -360 -243 -264 -209
rect 264 -243 360 -209
<< properties >>
string FIXED_BBOX -343 -226 343 226
<< end >>
