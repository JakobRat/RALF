magic
tech sky130A
magscale 1 2
timestamp 1702541237
<< checkpaint >>
rect -1556 -1997 1556 1997
<< nwell >>
rect -296 -737 296 737
<< pmos >>
rect -100 118 100 518
rect -100 -518 100 -118
<< pdiff >>
rect -158 506 -100 518
rect -158 130 -146 506
rect -112 130 -100 506
rect -158 118 -100 130
rect 100 506 158 518
rect 100 130 112 506
rect 146 130 158 506
rect 100 118 158 130
rect -158 -130 -100 -118
rect -158 -506 -146 -130
rect -112 -506 -100 -130
rect -158 -518 -100 -506
rect 100 -130 158 -118
rect 100 -506 112 -130
rect 146 -506 158 -130
rect 100 -518 158 -506
<< pdiffc >>
rect -146 130 -112 506
rect 112 130 146 506
rect -146 -506 -112 -130
rect 112 -506 146 -130
<< nsubdiff >>
rect -260 667 260 701
rect -260 -667 -226 667
rect 226 -667 260 667
rect -260 -701 -164 -667
rect 164 -701 260 -667
<< nsubdiffcont >>
rect -164 -701 164 -667
<< poly >>
rect -100 599 100 615
rect -100 565 -84 599
rect 84 565 100 599
rect -100 518 100 565
rect -100 71 100 118
rect -100 37 -84 71
rect 84 37 100 71
rect -100 21 100 37
rect -100 -37 100 -21
rect -100 -71 -84 -37
rect 84 -71 100 -37
rect -100 -118 100 -71
rect -100 -565 100 -518
rect -100 -599 -84 -565
rect 84 -599 100 -565
rect -100 -615 100 -599
<< polycont >>
rect -84 565 84 599
rect -84 37 84 71
rect -84 -71 84 -37
rect -84 -599 84 -565
<< locali >>
rect -260 667 260 701
rect -260 -667 -226 667
rect -100 565 -84 599
rect 84 565 100 599
rect -146 506 -112 522
rect -146 114 -112 130
rect 112 506 146 522
rect 112 114 146 130
rect -100 37 -84 71
rect 84 37 100 71
rect -100 -71 -84 -37
rect 84 -71 100 -37
rect -146 -130 -112 -114
rect -146 -522 -112 -506
rect 112 -130 146 -114
rect 112 -522 146 -506
rect -100 -599 -84 -565
rect 84 -599 100 -565
rect 226 -667 260 667
rect -260 -701 -164 -667
rect 164 -701 260 -667
<< properties >>
string FIXED_BBOX -243 -684 243 684
<< end >>
