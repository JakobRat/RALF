magic
tech sky130A
magscale 1 2
timestamp 1699959963
<< checkpaint >>
rect -357 1797 3013 4385
rect -1685 233 3013 1797
rect -1685 -325 2984 233
rect -1685 -1797 1685 -325
use XDL_XM3_XM4  XDL_XM3_XM4_0 ~/Documents/RALF/Magic/Devices
timestamp 1699959914
transform 1 0 1328 0 1 2588
box -425 -537 425 537
use XDP_XM1_XM2  XDP_XM1_XM2_0 ~/Documents/RALF/Magic/Devices
timestamp 1699959914
transform 1 0 1328 0 1 1772
box -425 -279 425 279
use XM5  XM5_0 ~/Documents/RALF/Magic/Devices
timestamp 1699959914
transform 1 0 1328 0 1 1214
box -396 -279 396 279
<< end >>
