** sch_path: /foss/designs/xschem/MillerOpAmp/OpAmp_tb.sch
**.subckt OpAmp_tb
V3 VDD GND 1.8
.save i(v3)
E1 Vp Vcmm vd GND 0.5
E2 Vn Vcmm vd GND -0.5
Vcmm Vcmm GND 0.9
.save i(vcmm)
Vd vd GND dc 0 ac 1
.save i(vd)
x1 VDD Vcmm Voutp Voutn Vp Vn GND OpAmp
C2 Voutn GND 50f m=1
C1 Voutp GND 50f m=1
**** begin user architecture code



* ngspice commands
.option savecurrents
.save all
.control
ac dec 1001 1 100Meg
let vod = V(Voutp)-V(Voutn)
meas ac gain max vod
let gain3dB = gain/sqrt(2)
meas ac BW TRIG at=1 TARG vod val=gain3dB fall=LAST
let GBW = BW*gain*1e-6
print GBW
print vodmax
plot vdb(vod) xlimit 1k 100Meg ylabel 'small signal gain'
let outd = 180/PI*cph(vod)
meas ac ftHz when vdb(vod)=1 fall=LAST
meas ac ph find outd when vdb(vod)=0 fall=LAST
let phm = ph+180
print phm
settype phase outd
plot outd xlimit 1k 100Meg ylabel 'phase'
dc Vd -0.02 0.02 1m
let vod = V(Voutp)-V(Voutn)
plot vod
op
write MillerOpAmp_tb.raw
.endc



 .lib /foss/pdks/sky130A/libs.tech/ngspice/sky130.lib.spice tt

**** end user architecture code
**.ends

* expanding   symbol:  /foss/designs/xschem/MillerOpAmp/OpAmp.sym # of pins=7
** sym_path: /foss/designs/xschem/MillerOpAmp/OpAmp.sym
** sch_path: /foss/designs/xschem/MillerOpAmp/OpAmp.sch
.subckt OpAmp VPWR Vcmm Vop Von Vp Vn VGND
*.opin Von
*.opin Vop
*.ipin Vcmm
*.ipin Vp
*.ipin Vn
*.iopin VPWR
*.iopin VGND
x1 VPWR Von Vcmmfb Vp Vn Vbias Vop VGND MillerOpAmp
x2 VPWR Vbias VGND Bias
x3 Vop VPWR Vcmm Vcmmfb Vbias VGND Von CMMFeedback
.ends


* expanding   symbol:  /foss/designs/xschem/MillerOpAmp/MillerOpAmp.sym # of pins=8
** sym_path: /foss/designs/xschem/MillerOpAmp/MillerOpAmp.sym
** sch_path: /foss/designs/xschem/MillerOpAmp/MillerOpAmp.sch
.subckt MillerOpAmp VPWR Von Vbias2 Vp Vn Vbias1 Vop VGND
*.opin Von
*.opin Vop
*.ipin Vbias2
*.ipin Vp
*.ipin Vn
*.ipin Vbias1
*.iopin VPWR
*.iopin VGND
XC1 Von1 Von sky130_fd_pr__cap_mim_m3_1 W=4 L=4 MF=1 m=1
XC2 Vop1 Vop sky130_fd_pr__cap_mim_m3_1 W=4 L=4 MF=1 m=1
x1 VPWR Vbias2 Von1 Vop1 Vp Vn Vbias1 VGND DiffAmp
x2 VPWR Von1 Von Vbias1 VGND CSAmp
x3 VPWR Vop1 Vop Vbias1 VGND CSAmp
.ends


* expanding   symbol:  /foss/designs/xschem/MillerOpAmp/Bias.sym # of pins=3
** sym_path: /foss/designs/xschem/MillerOpAmp/Bias.sym
** sch_path: /foss/designs/xschem/MillerOpAmp/Bias.sch
.subckt Bias Vdd Vbias Vss
*.opin Vbias
*.iopin Vss
*.iopin Vdd
XM6 Vbias Vbias Vss Vss sky130_fd_pr__nfet_01v8 L=2 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM2 VbiasP VbiasP Vdd Vdd sky130_fd_pr__pfet_01v8 L=2 W=1 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XR1 VbiasP net1 Vss sky130_fd_pr__res_xhigh_po_0p35 L=2 mult=1 m=1
XR2 net1 net2 Vss sky130_fd_pr__res_xhigh_po_0p35 L=2 mult=1 m=1
XR3 net2 net3 Vss sky130_fd_pr__res_xhigh_po_0p35 L=2 mult=1 m=1
XR4 net3 net4 Vss sky130_fd_pr__res_xhigh_po_0p35 L=2 mult=1 m=1
XR5 net4 Vbias Vss sky130_fd_pr__res_xhigh_po_0p35 L=2 mult=1 m=1
.ends


* expanding   symbol:  /foss/designs/xschem/MillerOpAmp/CMMFeedback.sym # of pins=7
** sym_path: /foss/designs/xschem/MillerOpAmp/CMMFeedback.sym
** sch_path: /foss/designs/xschem/MillerOpAmp/CMMFeedback.sch
.subckt CMMFeedback Vop Vdd Vcmm Vout Vbias Vss Von
*.ipin Vbias
*.opin Vout
*.ipin Vop
*.ipin Vcmm
*.ipin Von
*.iopin Vss
*.iopin Vdd
x2 Vdd net1 Vout net1 Vcmm VcmmOut Vbias Vss DiffAmp
XR6 Vop net2 Vss sky130_fd_pr__res_xhigh_po_0p35 L=2 mult=1 m=1
XR7 net2 net3 Vss sky130_fd_pr__res_xhigh_po_0p35 L=2 mult=1 m=1
XR8 net3 net4 Vss sky130_fd_pr__res_xhigh_po_0p35 L=2 mult=1 m=1
XR9 net4 net5 Vss sky130_fd_pr__res_xhigh_po_0p35 L=2 mult=1 m=1
XR10 net5 VcmmOut Vss sky130_fd_pr__res_xhigh_po_0p35 L=2 mult=1 m=1
XR11 Von net6 Vss sky130_fd_pr__res_xhigh_po_0p35 L=2 mult=1 m=1
XR12 net6 net7 Vss sky130_fd_pr__res_xhigh_po_0p35 L=2 mult=1 m=1
XR13 net7 net8 Vss sky130_fd_pr__res_xhigh_po_0p35 L=2 mult=1 m=1
XR14 net8 net9 Vss sky130_fd_pr__res_xhigh_po_0p35 L=2 mult=1 m=1
XR15 net9 VcmmOut Vss sky130_fd_pr__res_xhigh_po_0p35 L=2 mult=1 m=1
.ends


* expanding   symbol:  /foss/designs/xschem/MillerOpAmp/DiffAmp.sym # of pins=8
** sym_path: /foss/designs/xschem/MillerOpAmp/DiffAmp.sym
** sch_path: /foss/designs/xschem/MillerOpAmp/DiffAmp.sch
.subckt DiffAmp Vdd Vbias2 Von Vop Vp Vn Vbias1 Vss
*.iopin Vdd
*.iopin Vss
*.ipin Vp
*.ipin Vn
*.ipin Vbias1
*.ipin Vbias2
*.opin Vop
*.opin Von
XM1 Vop Vp Vmid Vss sky130_fd_pr__nfet_01v8 L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM2 Von Vn Vmid Vss sky130_fd_pr__nfet_01v8 L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM3 Vop Vbias2 Vdd Vdd sky130_fd_pr__pfet_01v8 L=1 W=2 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM4 Von Vbias2 Vdd Vdd sky130_fd_pr__pfet_01v8 L=1 W=2 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM5 Vmid Vbias1 Vss Vss sky130_fd_pr__nfet_01v8 L=2 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  /foss/designs/xschem/MillerOpAmp/CSAmp.sym # of pins=5
** sym_path: /foss/designs/xschem/MillerOpAmp/CSAmp.sym
** sch_path: /foss/designs/xschem/MillerOpAmp/CSAmp.sch
.subckt CSAmp Vdd Vi Vo Vbias1 Vss
*.ipin Vbias1
*.ipin Vi
*.iopin Vdd
*.iopin Vss
*.opin Vo
XM1 Vo Vi Vdd Vdd sky130_fd_pr__pfet_01v8 L=1 W=4 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM2 Vo Vbias1 Vss Vss sky130_fd_pr__nfet_01v8 L=2 W=12 nf=6 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
.ends

.GLOBAL GND
.GLOBAL VDD
.end
