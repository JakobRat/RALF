magic
tech sky130A
magscale 1 2
timestamp 1699960391
<< checkpaint >>
rect -1685 -1539 1685 1539
<< pwell >>
rect -425 -279 425 279
<< nmos >>
rect -229 -131 -29 69
rect 29 -131 229 69
<< ndiff >>
rect -287 57 -229 69
rect -287 -119 -275 57
rect -241 -119 -229 57
rect -287 -131 -229 -119
rect -29 57 29 69
rect -29 -119 -17 57
rect 17 -119 29 57
rect -29 -131 29 -119
rect 229 57 287 69
rect 229 -119 241 57
rect 275 -119 287 57
rect 229 -131 287 -119
<< ndiffc >>
rect -275 -119 -241 57
rect -17 -119 17 57
rect 241 -119 275 57
<< psubdiff >>
rect -389 209 389 243
rect -389 -209 -355 209
rect 355 -209 389 209
rect -389 -243 -293 -209
rect 293 -243 389 -209
<< psubdiffcont >>
rect -293 -243 293 -209
<< poly >>
rect -229 141 -29 157
rect -229 107 -213 141
rect -45 107 -29 141
rect -229 69 -29 107
rect 29 141 229 157
rect 29 107 45 141
rect 213 107 229 141
rect 29 69 229 107
rect -229 -157 -29 -131
rect 29 -157 229 -131
<< polycont >>
rect -213 107 -45 141
rect 45 107 213 141
<< locali >>
rect -389 209 389 243
rect -389 -209 -355 209
rect -229 107 -213 141
rect -45 107 -29 141
rect 29 107 45 141
rect 213 107 229 141
rect -275 57 -241 73
rect -275 -135 -241 -119
rect -17 57 17 73
rect -17 -135 17 -119
rect 241 57 275 73
rect 241 -135 275 -119
rect 355 -209 389 209
rect -389 -243 -293 -209
rect 293 -243 389 -209
<< properties >>
string FIXED_BBOX -372 -226 372 226
<< end >>
