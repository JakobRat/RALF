** sch_path: /home/jakob/Documents/RALF/Circuits/Examples/Latch/CCLatch_tb.sch
**.subckt CCLatch_tb
x1 VDD out outn in inn clk GND CCLatch
V1 VDD GND 1.8
.save i(v1)
V2 clk GND PULSE(0 1.8 50n 0.1n 0.1n 50ns 100ns 10)
.save i(v2)
V3 in GND PULSE(0 1.8 40ns 0.1n 0.1n 70ns 200ns 5)
.save i(v3)
E1 net1 GND in GND -1
V4 inn net1 1.8
.save i(v4)
**** begin user architecture code



* ngspice commands
.option savecurrents
.save all
.control
tran 10ns 1000ns
.endc



 .lib /home/jakob/pdks/sky130A/libs.tech/ngspice/sky130.lib.spice tt

**** end user architecture code
**.ends

* expanding   symbol:  /home/jakob/Documents/RALF/Circuits/Examples/Latch/CCLatch.sym # of pins=7
** sym_path: /home/jakob/Documents/RALF/Circuits/Examples/Latch/CCLatch.sym
** sch_path: /home/jakob/Documents/RALF/Circuits/Examples/Latch/CCLatch.sch
.subckt CCLatch Vdd out outn in inn clk Vss
*.iopin Vdd
*.iopin Vss
*.ipin in
*.ipin inn
*.ipin clk
*.opin outn
*.opin out
XM1 outn in Vmid Vss sky130_fd_pr__nfet_01v8 L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM2 out inn Vmid Vss sky130_fd_pr__nfet_01v8 L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM3 outn out Vdd Vdd sky130_fd_pr__pfet_01v8 L=1 W=2 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM4 out outn Vdd Vdd sky130_fd_pr__pfet_01v8 L=1 W=2 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM5 Vmid clk Vss Vss sky130_fd_pr__nfet_01v8 L=2 W=10 nf=5 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
.ends

.GLOBAL VDD
.GLOBAL GND
.end
