** sch_path: /home/jakob/Documents/AutomatedLayoutGeneration/Circuits/Buffer/Buffer.sch
**.subckt Buffer in out VPWR VGND
*.ipin in
*.opin out
*.iopin VPWR
*.iopin VGND
x1 VPWR in vo1 VGND inverter
x2 VPWR vo1 out VGND inverter
**.ends

* expanding   symbol:  /home/jakob/Documents/AutomatedLayoutGeneration/Circuits/Buffer/inverter.sym
*+ # of pins=4
** sym_path: /home/jakob/Documents/AutomatedLayoutGeneration/Circuits/Buffer/inverter.sym
** sch_path: /home/jakob/Documents/AutomatedLayoutGeneration/Circuits/Buffer/inverter.sch
.subckt inverter Vdd in out Vss
*.iopin Vdd
*.iopin Vss
*.ipin in
*.opin out
XM1 out in Vdd Vdd sky130_fd_pr__pfet_01v8 L=0.3 W='1 * 8 ' nf=8 ad='int((nf+1)/2) * W / nf * 0.29' as='int((nf+2)/2) * W / nf * 0.29'
+ pd='2*int((nf+1)/2) * (W / nf + 0.29)' ps='2*int((nf+2)/2) * (W / nf + 0.29)' nrd='0.29 / W ' nrs='0.29 / W '
+ sa=0 sb=0 sd=0 mult=1 m=1
XM2 out in Vss Vss sky130_fd_pr__nfet_01v8 L=0.3 W='1 * 8 ' nf=8 ad='int((nf+1)/2) * W / nf * 0.29' as='int((nf+2)/2) * W / nf * 0.29'
+ pd='2*int((nf+1)/2) * (W / nf + 0.29)' ps='2*int((nf+2)/2) * (W / nf + 0.29)' nrd='0.29 / W ' nrs='0.29 / W '
+ sa=0 sb=0 sd=0 mult=1 m=1
.ends

.end