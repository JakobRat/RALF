magic
tech sky130A
magscale 1 2
timestamp 1702977093
<< checkpaint >>
rect -1685 -1997 1685 1997
<< nwell >>
rect -425 -737 425 737
<< pmos >>
rect -229 118 -29 518
rect 29 118 229 518
rect -229 -518 -29 -118
rect 29 -518 229 -118
<< pdiff >>
rect -287 506 -229 518
rect -287 130 -275 506
rect -241 130 -229 506
rect -287 118 -229 130
rect -29 506 29 518
rect -29 130 -17 506
rect 17 130 29 506
rect -29 118 29 130
rect 229 506 287 518
rect 229 130 241 506
rect 275 130 287 506
rect 229 118 287 130
rect -287 -130 -229 -118
rect -287 -506 -275 -130
rect -241 -506 -229 -130
rect -287 -518 -229 -506
rect -29 -130 29 -118
rect -29 -506 -17 -130
rect 17 -506 29 -130
rect -29 -518 29 -506
rect 229 -130 287 -118
rect 229 -506 241 -130
rect 275 -506 287 -130
rect 229 -518 287 -506
<< pdiffc >>
rect -275 130 -241 506
rect -17 130 17 506
rect 241 130 275 506
rect -275 -506 -241 -130
rect -17 -506 17 -130
rect 241 -506 275 -130
<< nsubdiff >>
rect -389 667 389 701
rect -389 -667 -355 667
rect 355 -667 389 667
rect -389 -701 -293 -667
rect 293 -701 389 -667
<< nsubdiffcont >>
rect -293 -701 293 -667
<< poly >>
rect -229 599 -29 615
rect -229 565 -213 599
rect -45 565 -29 599
rect -229 518 -29 565
rect 29 599 229 615
rect 29 565 45 599
rect 213 565 229 599
rect 29 518 229 565
rect -229 71 -29 118
rect -229 37 -213 71
rect -45 37 -29 71
rect -229 21 -29 37
rect 29 71 229 118
rect 29 37 45 71
rect 213 37 229 71
rect 29 21 229 37
rect -229 -37 -29 -21
rect -229 -71 -213 -37
rect -45 -71 -29 -37
rect -229 -118 -29 -71
rect 29 -37 229 -21
rect 29 -71 45 -37
rect 213 -71 229 -37
rect 29 -118 229 -71
rect -229 -565 -29 -518
rect -229 -599 -213 -565
rect -45 -599 -29 -565
rect -229 -615 -29 -599
rect 29 -565 229 -518
rect 29 -599 45 -565
rect 213 -599 229 -565
rect 29 -615 229 -599
<< polycont >>
rect -213 565 -45 599
rect 45 565 213 599
rect -213 37 -45 71
rect 45 37 213 71
rect -213 -71 -45 -37
rect 45 -71 213 -37
rect -213 -599 -45 -565
rect 45 -599 213 -565
<< locali >>
rect -389 667 389 701
rect -389 -667 -355 667
rect -229 565 -213 599
rect -45 565 -29 599
rect 29 565 45 599
rect 213 565 229 599
rect -275 506 -241 522
rect -275 114 -241 130
rect -17 506 17 522
rect -17 114 17 130
rect 241 506 275 522
rect 241 114 275 130
rect -229 37 -213 71
rect -45 37 -29 71
rect 29 37 45 71
rect 213 37 229 71
rect -229 -71 -213 -37
rect -45 -71 -29 -37
rect 29 -71 45 -37
rect 213 -71 229 -37
rect -275 -130 -241 -114
rect -275 -522 -241 -506
rect -17 -130 17 -114
rect -17 -522 17 -506
rect 241 -130 275 -114
rect 241 -522 275 -506
rect -229 -599 -213 -565
rect -45 -599 -29 -565
rect 29 -599 45 -565
rect 213 -599 229 -565
rect 355 -667 389 667
rect -389 -701 -293 -667
rect 293 -701 389 -667
<< properties >>
string FIXED_BBOX -372 -684 372 684
<< end >>
