magic
tech sky130A
magscale 1 2
timestamp 1703087217
<< checkpaint >>
rect 617 2989 3695 3223
rect -233 2431 3695 2989
rect -545 1997 3695 2431
rect -1556 1556 3695 1997
rect -1997 -89 3695 1556
rect -1997 -681 3449 -89
rect -1997 -1556 1997 -681
rect -1556 -1997 1556 -1556
use XDL_XM3_XM4  XDL_XM3_XM4_0 ~/Documents/RALF/Magic/Devices
timestamp 1703087211
transform 0 -1 1452 1 0 875
box -296 -737 296 737
use XDP_XM1_XM2  XDP_XM1_XM2_0 ~/Documents/RALF/Magic/Devices
timestamp 1703087211
transform -1 0 1452 0 -1 1450
box -425 -279 425 279
use XM5  XM5_0 ~/Documents/RALF/Magic/Devices
timestamp 1703087211
transform 0 1 2156 -1 0 1567
box -396 -279 396 279
<< end >>
