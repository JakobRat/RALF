* expanding   symbol:
*+  /home/jakob/Documents/AutomatedLayoutGeneration/Circuits/Comparator/DiffAmp.sym # of pins=7
** sym_path: /home/jakob/Documents/AutomatedLayoutGeneration/Circuits/Comparator/DiffAmp.sym
** sch_path: /home/jakob/Documents/AutomatedLayoutGeneration/Circuits/Comparator/DiffAmp.sch
**.subckt DiffAmp clk VPWR outn outp inn inp VGND
*.iopin VPWR
*.iopin VGND
*.ipin clk
*.ipin inp
*.ipin inn
*.opin outn
*.opin outp
XM3 outn inp in_stage_net1 VGND sky130_fd_pr__nfet_01v8 L=0.3 W=8 nf=4 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM4 outp inn in_stage_net1 VGND sky130_fd_pr__nfet_01v8 L=0.3 W=8 nf=4 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM5 in_stage_net1 clk VGND VGND sky130_fd_pr__nfet_01v8 L=0.3 W=6 nf=6 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM2 outp clk VPWR VPWR sky130_fd_pr__pfet_01v8 L=0.3 W=3 nf=3 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM1 outn clk VPWR VPWR sky130_fd_pr__pfet_01v8 L=0.3 W=3 nf=3 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
**.ends
.end