magic
tech sky130A
magscale 1 2
timestamp 1701367482
<< checkpaint >>
rect -443 2673 3151 4081
rect -498 1797 3151 2673
rect -1685 1685 3151 1797
rect -1797 711 3151 1685
rect -1797 153 3061 711
rect -1797 -405 2814 153
rect -1797 -1685 1797 -405
rect -1685 -1797 1685 -1685
use XDL_XM3_XM4  XDL_XM3_XM4_0 ~/Documents/RALF/Magic/Devices
timestamp 1701367472
transform 0 1 1354 -1 0 2396
box -425 -537 425 537
use XDP_XM1_XM2  XDP_XM1_XM2_0 ~/Documents/RALF/Magic/Devices
timestamp 1701367472
transform 1 0 1376 0 1 1692
box -425 -279 425 279
use XM5  XM5_0 ~/Documents/RALF/Magic/Devices
timestamp 1701367472
transform -1 0 1158 0 -1 1134
box -396 -279 396 279
<< end >>
