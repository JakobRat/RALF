** sch_path:
*+ /home/jakob/Documents/AutomatedLayoutGeneration/Circuits/DiffAmp/TwoStageDiffAmp_flat.sch
**.subckt TwoStageDiffAmp_flat Vss Vn Vp Vout Vdd
*.iopin Vss
*.ipin Vn
*.ipin Vp
*.opin Vout
*.iopin Vdd
XR3 Vbias Vdd Vss sky130_fd_pr__res_xhigh_po_0p35 L=0.35 mult=1 m=1
XM4 Vbias Vbias Vss Vss sky130_fd_pr__nfet_01v8 L=0.3 W=0.84 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM1 Vo_p Vo_p Vdd VB1 sky130_fd_pr__pfet_01v8 L=0.3 W=0.84 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM2 Vo_n Vo_p Vdd VB1 sky130_fd_pr__pfet_01v8 L=0.3 W=0.84 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM3 Vo_p Vn Vmid Vss sky130_fd_pr__nfet_01v8 L=0.3 W=0.84 nf=5 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM5 Vo_n Vp Vmid Vss sky130_fd_pr__nfet_01v8 L=0.3 W=0.84 nf=5 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM6 Vmid Vbias Vss Vss sky130_fd_pr__nfet_01v8 L=0.3 W=0.84 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM7 Vout Vo_n Vdd Vdd sky130_fd_pr__pfet_01v8 L=0.3 W=0.84 nf=10 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XR4 Vss Vout Vss sky130_fd_pr__res_xhigh_po_0p35 L=20 mult=1 m=1
XC1 Vo_n Vout sky130_fd_pr__cap_mim_m3_1 W=2 L=2 MF=1 m=1
XC2 Vo_n Vout sky130_fd_pr__cap_mim_m3_1 W=2 L=2 MF=1 m=1
**.ends
.end