magic
tech sky130A
magscale 1 2
timestamp 1702720036
<< checkpaint >>
rect -1685 -1739 1685 1739
<< pwell >>
rect -425 -479 425 479
<< nmos >>
rect -229 -331 -29 269
rect 29 -331 229 269
<< ndiff >>
rect -287 257 -229 269
rect -287 -319 -275 257
rect -241 -319 -229 257
rect -287 -331 -229 -319
rect -29 257 29 269
rect -29 -319 -17 257
rect 17 -319 29 257
rect -29 -331 29 -319
rect 229 257 287 269
rect 229 -319 241 257
rect 275 -319 287 257
rect 229 -331 287 -319
<< ndiffc >>
rect -275 -319 -241 257
rect -17 -319 17 257
rect 241 -319 275 257
<< psubdiff >>
rect -389 409 389 443
rect -389 -409 -355 409
rect 355 -409 389 409
rect -389 -443 -293 -409
rect 293 -443 389 -409
<< psubdiffcont >>
rect -293 -443 293 -409
<< poly >>
rect -229 341 -29 357
rect -229 307 -213 341
rect -45 307 -29 341
rect -229 269 -29 307
rect 29 341 229 357
rect 29 307 45 341
rect 213 307 229 341
rect 29 269 229 307
rect -229 -357 -29 -331
rect 29 -357 229 -331
<< polycont >>
rect -213 307 -45 341
rect 45 307 213 341
<< locali >>
rect -389 409 389 443
rect -389 -409 -355 409
rect -229 307 -213 341
rect -45 307 -29 341
rect 29 307 45 341
rect 213 307 229 341
rect -275 257 -241 273
rect -275 -335 -241 -319
rect -17 257 17 273
rect -17 -335 17 -319
rect 241 257 275 273
rect 241 -335 275 -319
rect 355 -409 389 409
rect -389 -443 -293 -409
rect 293 -443 389 -409
<< properties >>
string FIXED_BBOX -372 -426 372 426
<< end >>
