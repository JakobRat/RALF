magic
tech sky130A
magscale 1 2
timestamp 1702058220
<< checkpaint >>
rect -179 2579 3191 3537
rect -445 2533 3191 2579
rect -445 1797 3517 2533
rect -1556 1739 3517 1797
rect -1685 -1061 3517 1739
rect -1685 -1739 1685 -1061
rect -1556 -1797 1556 -1739
use XCCP_XM3_XM4  XCCP_XM3_XM4_0 ~/Documents/RALF/Magic/Devices
timestamp 1702049922
transform 1 0 1961 0 1 736
box -296 -537 296 537
use XDP_XM1_XM2  XDP_XM1_XM2_0 ~/Documents/RALF/Magic/Devices
timestamp 1702049922
transform -1 0 1240 0 -1 840
box -425 -479 425 479
use XM5  XM5_0 ~/Documents/RALF/Magic/Devices
timestamp 1702049922
transform 1 0 1506 0 1 1798
box -425 -479 425 479
<< end >>
