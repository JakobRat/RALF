magic
tech sky130A
magscale 1 2
timestamp 1702067089
<< checkpaint >>
rect -1793 -2033 1793 2033
<< pwell >>
rect -533 -773 533 773
<< psubdiff >>
rect -497 703 497 737
rect -497 -703 -463 703
rect 463 -703 497 703
rect -497 -737 -401 -703
rect 401 -737 497 -703
<< psubdiffcont >>
rect -401 -737 401 -703
<< xpolycontact >>
rect -367 175 -297 607
rect -367 -607 -297 -175
rect -201 175 -131 607
rect -201 -607 -131 -175
rect -35 175 35 607
rect -35 -607 35 -175
rect 131 175 201 607
rect 131 -607 201 -175
rect 297 175 367 607
rect 297 -607 367 -175
<< xpolyres >>
rect -367 -175 -297 175
rect -201 -175 -131 175
rect -35 -175 35 175
rect 131 -175 201 175
rect 297 -175 367 175
<< locali >>
rect -417 -737 -401 -703
rect 401 -737 417 -703
<< res0p35 >>
rect -369 -177 -295 177
rect -203 -177 -129 177
rect -37 -177 37 177
rect 129 -177 203 177
rect 295 -177 369 177
<< properties >>
string FIXED_BBOX -480 -720 480 720
<< end >>
