magic
tech sky130A
magscale 1 2
timestamp 1702029109
<< checkpaint >>
rect 1438 3867 4550 4325
rect 1438 1997 5400 3867
rect -1556 1539 5400 1997
rect -1685 789 5400 1539
rect -1685 331 5342 789
rect -1685 -1539 1685 331
rect 2030 231 5342 331
rect -1556 -1997 1556 -1539
use XDL_XM3_XM4  XDL_XM3_XM4_0 ~/Documents/RALF/Magic/Devices
timestamp 1702029005
transform -1 0 2994 0 -1 2328
box -296 -737 296 737
use XDP_XM1_XM2  XDP_XM1_XM2_0 ~/Documents/RALF/Magic/Devices
timestamp 1702029005
transform -1 0 3715 0 -1 2328
box -425 -279 425 279
use XM5  XM5_0 ~/Documents/RALF/Magic/Devices
timestamp 1702029005
transform -1 0 3686 0 -1 1770
box -396 -279 396 279
<< end >>
