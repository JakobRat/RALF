magic
tech sky130A
magscale 1 2
timestamp 1691681432
<< metal1 >>
rect 4808 11284 4872 11290
rect 4808 11232 4814 11284
rect 4866 11232 4872 11284
rect 4808 11226 4872 11232
rect 5270 11224 5328 11230
rect 5322 11172 5328 11224
rect 5270 11166 5328 11172
rect 5270 11106 5328 11112
rect 5322 11054 5328 11106
rect 4808 11048 4872 11054
rect 5270 11048 5328 11054
rect 4808 10996 4814 11048
rect 4866 10996 4872 11048
rect 4808 10990 4872 10996
rect 5270 10988 5328 10994
rect 5322 10936 5328 10988
rect 5270 10930 5328 10936
rect 5270 10870 5328 10876
rect 5322 10818 5328 10870
rect 4808 10812 4872 10818
rect 5270 10812 5328 10818
rect 4808 10760 4814 10812
rect 4866 10760 4872 10812
rect 4808 10754 4872 10760
rect 4808 10478 4872 10484
rect 4808 10426 4814 10478
rect 4866 10426 4872 10478
rect 4808 10420 4872 10426
rect 5270 10418 5328 10424
rect 5322 10366 5328 10418
rect 5270 10360 5328 10366
rect 5270 10300 5328 10306
rect 5322 10248 5328 10300
rect 4808 10242 4872 10248
rect 5270 10242 5328 10248
rect 4808 10190 4814 10242
rect 4866 10190 4872 10242
rect 4808 10184 4872 10190
rect 5270 10182 5328 10188
rect 5322 10130 5328 10182
rect 5270 10124 5328 10130
rect 5270 10064 5328 10070
rect 5322 10012 5328 10064
rect 4808 10006 4872 10012
rect 5270 10006 5328 10012
rect 4808 9954 4814 10006
rect 4866 9954 4872 10006
rect 4808 9948 4872 9954
rect 4808 9672 4872 9678
rect 4808 9620 4814 9672
rect 4866 9620 4872 9672
rect 4808 9614 4872 9620
rect 5270 9612 5328 9618
rect 5322 9560 5328 9612
rect 5270 9554 5328 9560
rect 5270 9494 5328 9500
rect 5322 9442 5328 9494
rect 4808 9436 4872 9442
rect 5270 9436 5328 9442
rect 4808 9384 4814 9436
rect 4866 9384 4872 9436
rect 4808 9378 4872 9384
rect 5270 9376 5328 9382
rect 5322 9324 5328 9376
rect 5270 9318 5328 9324
rect 5270 9258 5328 9264
rect 5322 9206 5328 9258
rect 4808 9200 4872 9206
rect 5270 9200 5328 9206
rect 4808 9148 4814 9200
rect 4866 9148 4872 9200
rect 4808 9142 4872 9148
rect 4804 8866 4868 8872
rect 4804 8814 4810 8866
rect 4862 8814 4868 8866
rect 4804 8808 4868 8814
rect 5268 8806 5332 8812
rect 5268 8754 5274 8806
rect 5326 8754 5332 8806
rect 5268 8748 5332 8754
rect 5268 8688 5332 8694
rect 5268 8636 5274 8688
rect 5326 8636 5332 8688
rect 4804 8630 4868 8636
rect 5268 8630 5332 8636
rect 4804 8578 4810 8630
rect 4862 8578 4868 8630
rect 4804 8572 4868 8578
rect 5268 8570 5332 8576
rect 5268 8518 5274 8570
rect 5326 8518 5332 8570
rect 5268 8512 5332 8518
rect 5268 8452 5332 8458
rect 5268 8400 5274 8452
rect 5326 8400 5332 8452
rect 4804 8394 4868 8400
rect 5268 8394 5332 8400
rect 4804 8342 4810 8394
rect 4862 8342 4868 8394
rect 4804 8336 4868 8342
rect 4566 8060 4630 8066
rect 4566 8008 4572 8060
rect 4624 8008 4630 8060
rect 4566 8002 4630 8008
rect 5030 8000 5094 8006
rect 5030 7948 5036 8000
rect 5088 7948 5094 8000
rect 5030 7942 5094 7948
rect 5030 7882 5094 7888
rect 5030 7830 5036 7882
rect 5088 7830 5094 7882
rect 4566 7824 4630 7830
rect 5030 7824 5094 7830
rect 4566 7772 4572 7824
rect 4624 7772 4630 7824
rect 4566 7766 4630 7772
rect 5030 7764 5094 7770
rect 5030 7712 5036 7764
rect 5088 7712 5094 7764
rect 5030 7706 5094 7712
rect 5030 7646 5094 7652
rect 5030 7594 5036 7646
rect 5088 7594 5094 7646
rect 4566 7588 4630 7594
rect 5030 7588 5094 7594
rect 4566 7536 4572 7588
rect 4624 7536 4630 7588
rect 4566 7530 4630 7536
rect 4566 7254 4630 7260
rect 4566 7202 4572 7254
rect 4624 7202 4630 7254
rect 4566 7196 4630 7202
rect 5030 7194 5094 7200
rect 5030 7142 5036 7194
rect 5088 7142 5094 7194
rect 5030 7136 5094 7142
rect 5030 7076 5094 7082
rect 5030 7024 5036 7076
rect 5088 7024 5094 7076
rect 4566 7018 4630 7024
rect 5030 7018 5094 7024
rect 4566 6966 4572 7018
rect 4624 6966 4630 7018
rect 4566 6960 4630 6966
rect 5030 6958 5094 6964
rect 5030 6906 5036 6958
rect 5088 6906 5094 6958
rect 5030 6900 5094 6906
rect 5030 6840 5094 6846
rect 5030 6788 5036 6840
rect 5088 6788 5094 6840
rect 4566 6782 4630 6788
rect 5030 6782 5094 6788
rect 4566 6730 4572 6782
rect 4624 6730 4630 6782
rect 4566 6724 4630 6730
rect 4566 6448 4630 6454
rect 4566 6396 4572 6448
rect 4624 6396 4630 6448
rect 4566 6390 4630 6396
rect 5030 6388 5094 6394
rect 5030 6336 5036 6388
rect 5088 6336 5094 6388
rect 5030 6330 5094 6336
rect 5030 6270 5094 6276
rect 5030 6218 5036 6270
rect 5088 6218 5094 6270
rect 4566 6212 4630 6218
rect 5030 6212 5094 6218
rect 4566 6160 4572 6212
rect 4624 6160 4630 6212
rect 4566 6154 4630 6160
rect 5030 6152 5094 6158
rect 5030 6100 5036 6152
rect 5088 6100 5094 6152
rect 5030 6094 5094 6100
rect 5030 6034 5094 6040
rect 5030 5982 5036 6034
rect 5088 5982 5094 6034
rect 4566 5976 4630 5982
rect 5030 5976 5094 5982
rect 4566 5924 4572 5976
rect 4624 5924 4630 5976
rect 4566 5918 4630 5924
rect 4570 5642 4634 5648
rect 4570 5590 4576 5642
rect 4628 5590 4634 5642
rect 4570 5584 4634 5590
rect 5032 5582 5090 5588
rect 5084 5530 5090 5582
rect 5032 5524 5090 5530
rect 5032 5464 5090 5470
rect 5084 5412 5090 5464
rect 4570 5406 4634 5412
rect 5032 5406 5090 5412
rect 4570 5354 4576 5406
rect 4628 5354 4634 5406
rect 4570 5348 4634 5354
rect 5032 5346 5090 5352
rect 5084 5294 5090 5346
rect 5032 5288 5090 5294
rect 5032 5228 5090 5234
rect 5084 5176 5090 5228
rect 4570 5170 4634 5176
rect 5032 5170 5090 5176
rect 4570 5118 4576 5170
rect 4628 5118 4634 5170
rect 4570 5112 4634 5118
rect 4570 4836 4634 4842
rect 4570 4784 4576 4836
rect 4628 4784 4634 4836
rect 4570 4778 4634 4784
rect 5032 4776 5090 4782
rect 5084 4724 5090 4776
rect 5032 4718 5090 4724
rect 5032 4658 5090 4664
rect 5084 4606 5090 4658
rect 4570 4600 4634 4606
rect 5032 4600 5090 4606
rect 4570 4548 4576 4600
rect 4628 4548 4634 4600
rect 4570 4542 4634 4548
rect 5032 4540 5090 4546
rect 5084 4488 5090 4540
rect 5032 4482 5090 4488
rect 5032 4422 5090 4428
rect 5084 4370 5090 4422
rect 4570 4364 4634 4370
rect 5032 4364 5090 4370
rect 4570 4312 4576 4364
rect 4628 4312 4634 4364
rect 4570 4306 4634 4312
rect 4566 4030 4630 4036
rect 4566 3978 4572 4030
rect 4624 3978 4630 4030
rect 4566 3972 4630 3978
rect 5030 3970 5094 3976
rect 5030 3918 5036 3970
rect 5088 3918 5094 3970
rect 5030 3912 5094 3918
rect 5030 3852 5094 3858
rect 5030 3800 5036 3852
rect 5088 3800 5094 3852
rect 4566 3794 4630 3800
rect 5030 3794 5094 3800
rect 4566 3742 4572 3794
rect 4624 3742 4630 3794
rect 4566 3736 4630 3742
rect 5030 3734 5094 3740
rect 5030 3682 5036 3734
rect 5088 3682 5094 3734
rect 5030 3676 5094 3682
rect 5030 3616 5094 3622
rect 5030 3564 5036 3616
rect 5088 3564 5094 3616
rect 4566 3558 4630 3564
rect 5030 3558 5094 3564
rect 4566 3506 4572 3558
rect 4624 3506 4630 3558
rect 4566 3500 4630 3506
<< via1 >>
rect 4814 11232 4866 11284
rect 5270 11172 5322 11224
rect 5270 11054 5322 11106
rect 4814 10996 4866 11048
rect 5270 10936 5322 10988
rect 5270 10818 5322 10870
rect 4814 10760 4866 10812
rect 4814 10426 4866 10478
rect 5270 10366 5322 10418
rect 5270 10248 5322 10300
rect 4814 10190 4866 10242
rect 5270 10130 5322 10182
rect 5270 10012 5322 10064
rect 4814 9954 4866 10006
rect 4814 9620 4866 9672
rect 5270 9560 5322 9612
rect 5270 9442 5322 9494
rect 4814 9384 4866 9436
rect 5270 9324 5322 9376
rect 5270 9206 5322 9258
rect 4814 9148 4866 9200
rect 4810 8814 4862 8866
rect 5274 8754 5326 8806
rect 5274 8636 5326 8688
rect 4810 8578 4862 8630
rect 5274 8518 5326 8570
rect 5274 8400 5326 8452
rect 4810 8342 4862 8394
rect 4572 8008 4624 8060
rect 5036 7948 5088 8000
rect 5036 7830 5088 7882
rect 4572 7772 4624 7824
rect 5036 7712 5088 7764
rect 5036 7594 5088 7646
rect 4572 7536 4624 7588
rect 4572 7202 4624 7254
rect 5036 7142 5088 7194
rect 5036 7024 5088 7076
rect 4572 6966 4624 7018
rect 5036 6906 5088 6958
rect 5036 6788 5088 6840
rect 4572 6730 4624 6782
rect 4572 6396 4624 6448
rect 5036 6336 5088 6388
rect 5036 6218 5088 6270
rect 4572 6160 4624 6212
rect 5036 6100 5088 6152
rect 5036 5982 5088 6034
rect 4572 5924 4624 5976
rect 4576 5590 4628 5642
rect 5032 5530 5084 5582
rect 5032 5412 5084 5464
rect 4576 5354 4628 5406
rect 5032 5294 5084 5346
rect 5032 5176 5084 5228
rect 4576 5118 4628 5170
rect 4576 4784 4628 4836
rect 5032 4724 5084 4776
rect 5032 4606 5084 4658
rect 4576 4548 4628 4600
rect 5032 4488 5084 4540
rect 5032 4370 5084 4422
rect 4576 4312 4628 4364
rect 4572 3978 4624 4030
rect 5036 3918 5088 3970
rect 5036 3800 5088 3852
rect 4572 3742 4624 3794
rect 5036 3682 5088 3734
rect 5036 3564 5088 3616
rect 4572 3506 4624 3558
<< metal2 >>
rect 4808 11284 4872 11295
rect 4808 11255 4814 11284
rect 4718 11246 4814 11255
rect 4718 11190 4726 11246
rect 4782 11232 4814 11246
rect 4866 11232 4872 11284
rect 4782 11221 4872 11232
rect 5222 11254 5296 11255
rect 5222 11246 5340 11254
rect 4782 11190 4840 11221
rect 4718 11181 4840 11190
rect 5222 11190 5230 11246
rect 5286 11224 5340 11246
rect 5222 11172 5270 11190
rect 5322 11172 5340 11224
rect 5222 11144 5340 11172
rect 5222 11088 5230 11144
rect 5286 11106 5340 11144
rect 4808 11051 4872 11059
rect 4718 11048 4872 11051
rect 4718 11042 4814 11048
rect 4718 10986 4726 11042
rect 4782 10996 4814 11042
rect 4866 10996 4872 11048
rect 4782 10986 4872 10996
rect 4718 10985 4872 10986
rect 5222 11054 5270 11088
rect 5322 11054 5340 11106
rect 5222 10988 5340 11054
rect 4718 10977 4840 10985
rect 5222 10940 5270 10988
rect 5222 10884 5230 10940
rect 5322 10936 5340 10988
rect 5286 10884 5340 10936
rect 5222 10870 5340 10884
rect 5222 10847 5270 10870
rect 3962 10838 4840 10847
rect 3962 10782 3970 10838
rect 4026 10782 4726 10838
rect 4782 10823 4840 10838
rect 4970 10838 5270 10847
rect 4782 10812 4872 10823
rect 4782 10782 4814 10812
rect 3962 10773 4814 10782
rect 4808 10760 4814 10773
rect 4866 10760 4872 10812
rect 4970 10782 4978 10838
rect 5034 10782 5230 10838
rect 5322 10818 5340 10870
rect 5286 10782 5340 10818
rect 4970 10773 5340 10782
rect 5222 10772 5340 10773
rect 4808 10749 4872 10760
rect 4808 10478 4872 10489
rect 4808 10439 4814 10478
rect 4718 10430 4814 10439
rect 4718 10374 4726 10430
rect 4782 10426 4814 10430
rect 4866 10439 4872 10478
rect 4866 10430 5042 10439
rect 5222 10438 5296 10439
rect 4866 10426 4978 10430
rect 4782 10374 4978 10426
rect 5034 10374 5042 10430
rect 4718 10365 5042 10374
rect 5220 10430 5338 10438
rect 5220 10374 5230 10430
rect 5286 10418 5338 10430
rect 5220 10366 5270 10374
rect 5322 10366 5338 10418
rect 5220 10328 5338 10366
rect 5220 10272 5230 10328
rect 5286 10300 5338 10328
rect 4808 10242 4872 10253
rect 4808 10235 4814 10242
rect 4718 10226 4814 10235
rect 4718 10170 4726 10226
rect 4782 10190 4814 10226
rect 4866 10190 4872 10242
rect 4782 10179 4872 10190
rect 5220 10248 5270 10272
rect 5322 10248 5338 10300
rect 5220 10226 5338 10248
rect 4782 10170 4840 10179
rect 4718 10161 4840 10170
rect 5220 10170 5230 10226
rect 5286 10182 5338 10226
rect 5220 10130 5270 10170
rect 5322 10130 5338 10182
rect 5220 10064 5338 10130
rect 5220 10031 5270 10064
rect 4466 10022 4840 10031
rect 4466 9966 4474 10022
rect 4530 9966 4726 10022
rect 4782 10017 4840 10022
rect 4970 10022 5270 10031
rect 4782 10006 4872 10017
rect 4782 9966 4814 10006
rect 4466 9957 4814 9966
rect 4808 9954 4814 9957
rect 4866 9954 4872 10006
rect 4970 9966 4978 10022
rect 5034 9966 5230 10022
rect 5322 10012 5338 10064
rect 5286 9966 5338 10012
rect 4970 9960 5338 9966
rect 4970 9957 5296 9960
rect 4808 9943 4872 9954
rect 4718 9716 5042 9725
rect 4718 9660 4726 9716
rect 4782 9672 4978 9716
rect 4782 9660 4814 9672
rect 4718 9651 4814 9660
rect 4808 9620 4814 9651
rect 4866 9660 4978 9672
rect 5034 9660 5042 9716
rect 4866 9651 5042 9660
rect 4866 9620 4872 9651
rect 4808 9609 4872 9620
rect 5214 9614 5332 9644
rect 5214 9558 5230 9614
rect 5286 9612 5332 9614
rect 5322 9560 5332 9612
rect 5286 9558 5332 9560
rect 5214 9512 5332 9558
rect 5214 9456 5230 9512
rect 5286 9494 5332 9512
rect 4808 9436 4872 9447
rect 4808 9419 4814 9436
rect 4718 9410 4814 9419
rect 4718 9354 4726 9410
rect 4782 9384 4814 9410
rect 4866 9384 4872 9436
rect 4782 9373 4872 9384
rect 5214 9442 5270 9456
rect 5322 9442 5332 9494
rect 5214 9410 5332 9442
rect 4782 9354 4840 9373
rect 4718 9345 4840 9354
rect 5214 9354 5230 9410
rect 5286 9376 5332 9410
rect 5214 9324 5270 9354
rect 5322 9324 5332 9376
rect 5214 9308 5332 9324
rect 5214 9252 5230 9308
rect 5286 9258 5332 9308
rect 4718 9206 5042 9215
rect 4718 9150 4726 9206
rect 4782 9200 4978 9206
rect 4782 9150 4814 9200
rect 4718 9148 4814 9150
rect 4866 9150 4978 9200
rect 5034 9150 5042 9206
rect 5214 9206 5270 9252
rect 5322 9206 5332 9258
rect 5214 9166 5332 9206
rect 4866 9148 5042 9150
rect 4718 9141 5042 9148
rect 4808 9137 4872 9141
rect 4466 8900 4838 8909
rect 4466 8844 4474 8900
rect 4530 8844 4726 8900
rect 4782 8877 4838 8900
rect 4782 8866 4868 8877
rect 4782 8844 4810 8866
rect 4466 8835 4810 8844
rect 4804 8814 4810 8835
rect 4862 8814 4868 8866
rect 4804 8803 4868 8814
rect 5220 8807 5338 8852
rect 4970 8806 5338 8807
rect 4970 8798 5274 8806
rect 4970 8742 4978 8798
rect 5034 8754 5274 8798
rect 5326 8754 5338 8806
rect 5034 8742 5338 8754
rect 4970 8733 5338 8742
rect 5220 8705 5338 8733
rect 4970 8696 5338 8705
rect 4804 8630 4868 8641
rect 4970 8640 4978 8696
rect 5034 8688 5338 8696
rect 5034 8640 5274 8688
rect 4970 8636 5274 8640
rect 5326 8636 5338 8688
rect 4970 8631 5338 8636
rect 4804 8603 4810 8630
rect 4718 8594 4810 8603
rect 4718 8538 4726 8594
rect 4782 8578 4810 8594
rect 4862 8578 4868 8630
rect 5220 8603 5338 8631
rect 4782 8567 4868 8578
rect 4970 8594 5338 8603
rect 4782 8538 4838 8567
rect 4718 8529 4838 8538
rect 4970 8538 4978 8594
rect 5034 8570 5338 8594
rect 5034 8538 5274 8570
rect 4970 8529 5274 8538
rect 5220 8518 5274 8529
rect 5326 8518 5338 8570
rect 5220 8501 5338 8518
rect 4970 8492 5338 8501
rect 4970 8436 4978 8492
rect 5034 8452 5338 8492
rect 5034 8436 5274 8452
rect 4970 8427 5274 8436
rect 4804 8399 4868 8405
rect 4214 8394 4868 8399
rect 4214 8390 4810 8394
rect 4214 8334 4222 8390
rect 4278 8334 4726 8390
rect 4782 8342 4810 8390
rect 4862 8342 4868 8394
rect 5220 8400 5274 8427
rect 5326 8400 5338 8452
rect 5220 8374 5338 8400
rect 4782 8334 4868 8342
rect 4214 8331 4868 8334
rect 4214 8325 4838 8331
rect 4718 8186 5042 8195
rect 4718 8130 4726 8186
rect 4782 8130 4978 8186
rect 5034 8130 5042 8186
rect 4718 8121 5042 8130
rect 4466 8084 4790 8093
rect 4466 8028 4474 8084
rect 4530 8060 4726 8084
rect 4530 8028 4572 8060
rect 4466 8019 4572 8028
rect 4566 8008 4572 8019
rect 4624 8028 4726 8060
rect 4782 8028 4790 8084
rect 4624 8019 4790 8028
rect 4624 8008 4630 8019
rect 4566 7997 4630 8008
rect 4986 8000 5104 8026
rect 4986 7991 5036 8000
rect 4970 7982 5036 7991
rect 4970 7926 4978 7982
rect 5034 7948 5036 7982
rect 5088 7991 5104 8000
rect 5088 7982 5294 7991
rect 5088 7948 5230 7982
rect 5034 7926 5230 7948
rect 5286 7926 5294 7982
rect 4970 7917 5294 7926
rect 4986 7889 5104 7917
rect 4970 7882 5104 7889
rect 4970 7880 5036 7882
rect 4566 7824 4630 7835
rect 4566 7787 4572 7824
rect 4466 7778 4572 7787
rect 4466 7722 4474 7778
rect 4530 7772 4572 7778
rect 4624 7772 4630 7824
rect 4970 7824 4978 7880
rect 5034 7830 5036 7880
rect 5088 7830 5104 7882
rect 5034 7824 5104 7830
rect 4970 7815 5104 7824
rect 4986 7787 5104 7815
rect 4530 7761 4630 7772
rect 4970 7778 5104 7787
rect 4530 7722 4598 7761
rect 4466 7713 4598 7722
rect 4970 7722 4978 7778
rect 5034 7764 5104 7778
rect 5034 7722 5036 7764
rect 4970 7713 5036 7722
rect 4986 7712 5036 7713
rect 5088 7712 5104 7764
rect 4986 7685 5104 7712
rect 4718 7676 5104 7685
rect 4718 7620 4726 7676
rect 4782 7620 4978 7676
rect 5034 7646 5104 7676
rect 5034 7620 5036 7646
rect 4718 7611 5036 7620
rect 4566 7588 4630 7599
rect 4566 7583 4572 7588
rect 4466 7574 4572 7583
rect 4466 7518 4474 7574
rect 4530 7536 4572 7574
rect 4624 7536 4630 7588
rect 4986 7594 5036 7611
rect 5088 7594 5104 7646
rect 4986 7548 5104 7594
rect 4530 7525 4630 7536
rect 4530 7518 4598 7525
rect 4466 7509 4598 7518
rect 4466 7268 4790 7277
rect 4466 7212 4474 7268
rect 4530 7254 4726 7268
rect 4530 7212 4572 7254
rect 4466 7203 4572 7212
rect 4566 7202 4572 7203
rect 4624 7212 4726 7254
rect 4782 7212 4790 7268
rect 4624 7203 4790 7212
rect 4624 7202 4630 7203
rect 4566 7191 4630 7202
rect 4980 7194 5098 7230
rect 4980 7175 5036 7194
rect 4970 7166 5036 7175
rect 4970 7110 4978 7166
rect 5034 7142 5036 7166
rect 5088 7142 5098 7194
rect 5034 7110 5098 7142
rect 4970 7101 5098 7110
rect 4980 7076 5098 7101
rect 4980 7073 5036 7076
rect 4466 7064 4598 7073
rect 4466 7008 4474 7064
rect 4530 7029 4598 7064
rect 4970 7064 5036 7073
rect 4530 7018 4630 7029
rect 4530 7008 4572 7018
rect 4466 6999 4572 7008
rect 4566 6966 4572 6999
rect 4624 6966 4630 7018
rect 4970 7008 4978 7064
rect 5034 7024 5036 7064
rect 5088 7024 5098 7076
rect 5034 7008 5098 7024
rect 4970 6999 5098 7008
rect 4980 6971 5098 6999
rect 4566 6955 4630 6966
rect 4970 6962 5098 6971
rect 4970 6906 4978 6962
rect 5034 6958 5098 6962
rect 5034 6906 5036 6958
rect 5088 6906 5098 6958
rect 4970 6897 5098 6906
rect 4980 6869 5098 6897
rect 4970 6860 5098 6869
rect 4970 6804 4978 6860
rect 5034 6840 5098 6860
rect 5034 6804 5036 6840
rect 4970 6795 5036 6804
rect 4566 6782 4630 6793
rect 4566 6767 4572 6782
rect 4466 6758 4572 6767
rect 4466 6702 4474 6758
rect 4530 6730 4572 6758
rect 4624 6730 4630 6782
rect 4980 6788 5036 6795
rect 5088 6788 5098 6840
rect 4980 6752 5098 6788
rect 4530 6719 4630 6730
rect 4530 6702 4598 6719
rect 4466 6693 4598 6702
rect 4214 6554 4790 6563
rect 4214 6498 4222 6554
rect 4278 6498 4726 6554
rect 4782 6498 4790 6554
rect 4214 6489 4790 6498
rect 3962 6459 4598 6461
rect 3962 6452 4630 6459
rect 3962 6396 3970 6452
rect 4026 6448 4630 6452
rect 4026 6396 4572 6448
rect 4624 6396 4630 6448
rect 3962 6387 4630 6396
rect 4566 6385 4630 6387
rect 5014 6388 5132 6444
rect 5014 6359 5036 6388
rect 4718 6350 5036 6359
rect 4718 6294 4726 6350
rect 4782 6336 5036 6350
rect 5088 6359 5132 6388
rect 5088 6350 5294 6359
rect 5088 6336 5230 6350
rect 4782 6294 5230 6336
rect 5286 6294 5294 6350
rect 4718 6285 5294 6294
rect 5014 6270 5132 6285
rect 3962 6248 4598 6257
rect 3962 6192 3970 6248
rect 4026 6192 4222 6248
rect 4278 6223 4598 6248
rect 4278 6212 4630 6223
rect 4278 6192 4572 6212
rect 3962 6183 4572 6192
rect 4566 6160 4572 6183
rect 4624 6160 4630 6212
rect 4566 6149 4630 6160
rect 5014 6218 5036 6270
rect 5088 6257 5132 6270
rect 5088 6248 5294 6257
rect 5088 6218 5230 6248
rect 5014 6192 5230 6218
rect 5286 6192 5294 6248
rect 5014 6183 5294 6192
rect 5014 6155 5132 6183
rect 5014 6152 5294 6155
rect 5014 6100 5036 6152
rect 5088 6146 5294 6152
rect 5088 6100 5230 6146
rect 5014 6090 5230 6100
rect 5286 6090 5294 6146
rect 5014 6081 5294 6090
rect 5014 6053 5132 6081
rect 5014 6044 5294 6053
rect 5014 6034 5230 6044
rect 4566 5976 4630 5987
rect 4566 5951 4572 5976
rect 4214 5942 4572 5951
rect 4214 5886 4222 5942
rect 4278 5924 4572 5942
rect 4624 5951 4630 5976
rect 5014 5982 5036 6034
rect 5088 5988 5230 6034
rect 5286 5988 5294 6044
rect 5088 5982 5294 5988
rect 5014 5979 5294 5982
rect 5014 5966 5132 5979
rect 4624 5942 4790 5951
rect 4624 5924 4726 5942
rect 4278 5886 4726 5924
rect 4782 5886 4790 5942
rect 4214 5877 4790 5886
rect 4718 5840 5294 5849
rect 4718 5784 4726 5840
rect 4782 5784 5230 5840
rect 5286 5784 5294 5840
rect 4718 5775 5294 5784
rect 4570 5645 4634 5653
rect 4466 5642 4634 5645
rect 4466 5636 4576 5642
rect 4466 5580 4474 5636
rect 4530 5590 4576 5636
rect 4628 5590 4634 5642
rect 4530 5580 4634 5590
rect 4466 5579 4634 5580
rect 4974 5582 5092 5620
rect 4466 5571 4602 5579
rect 4974 5543 5032 5582
rect 4970 5534 5032 5543
rect 4970 5478 4978 5534
rect 5084 5530 5092 5582
rect 5034 5478 5092 5530
rect 4970 5469 5092 5478
rect 4974 5464 5092 5469
rect 4974 5441 5032 5464
rect 4466 5432 4602 5441
rect 4466 5376 4474 5432
rect 4530 5417 4602 5432
rect 4970 5432 5032 5441
rect 4530 5406 4634 5417
rect 4530 5376 4576 5406
rect 4466 5367 4576 5376
rect 4570 5354 4576 5367
rect 4628 5354 4634 5406
rect 4970 5376 4978 5432
rect 5084 5412 5092 5464
rect 5034 5376 5092 5412
rect 4970 5367 5092 5376
rect 4570 5343 4634 5354
rect 4974 5346 5092 5367
rect 4974 5339 5032 5346
rect 4970 5330 5032 5339
rect 4970 5274 4978 5330
rect 5084 5294 5092 5346
rect 5034 5274 5092 5294
rect 4970 5265 5092 5274
rect 4974 5237 5092 5265
rect 4718 5228 5092 5237
rect 4570 5170 4634 5181
rect 4570 5135 4576 5170
rect 4466 5126 4576 5135
rect 4466 5070 4474 5126
rect 4530 5118 4576 5126
rect 4628 5118 4634 5170
rect 4718 5172 4726 5228
rect 4782 5172 4978 5228
rect 5084 5176 5092 5228
rect 5034 5172 5092 5176
rect 4718 5163 5092 5172
rect 4974 5142 5092 5163
rect 4530 5107 4634 5118
rect 4530 5070 4602 5107
rect 4466 5061 4602 5070
rect 4570 4836 4634 4847
rect 4570 4829 4576 4836
rect 4466 4820 4576 4829
rect 4466 4764 4474 4820
rect 4530 4784 4576 4820
rect 4628 4829 4634 4836
rect 4628 4820 4790 4829
rect 4628 4784 4726 4820
rect 4530 4764 4726 4784
rect 4782 4764 4790 4820
rect 4466 4755 4790 4764
rect 4970 4820 5294 4829
rect 4970 4764 4978 4820
rect 5034 4776 5230 4820
rect 5084 4764 5230 4776
rect 5286 4764 5294 4820
rect 4970 4755 5032 4764
rect 4974 4724 5032 4755
rect 5084 4755 5294 4764
rect 5084 4724 5092 4755
rect 4974 4658 5092 4724
rect 4974 4625 5032 4658
rect 4466 4616 4602 4625
rect 4466 4560 4474 4616
rect 4530 4611 4602 4616
rect 4970 4616 5032 4625
rect 4530 4600 4634 4611
rect 4530 4560 4576 4600
rect 4466 4551 4576 4560
rect 4570 4548 4576 4551
rect 4628 4548 4634 4600
rect 4970 4560 4978 4616
rect 5084 4606 5092 4658
rect 5034 4560 5092 4606
rect 4970 4551 5092 4560
rect 4570 4537 4634 4548
rect 4974 4540 5092 4551
rect 4974 4523 5032 4540
rect 4970 4514 5032 4523
rect 4970 4458 4978 4514
rect 5084 4488 5092 4540
rect 5034 4458 5092 4488
rect 4970 4449 5092 4458
rect 4974 4422 5092 4449
rect 4974 4421 5032 4422
rect 4466 4412 4602 4421
rect 4466 4356 4474 4412
rect 4530 4375 4602 4412
rect 4970 4412 5032 4421
rect 4530 4364 4634 4375
rect 4530 4356 4576 4364
rect 4466 4347 4576 4356
rect 4570 4312 4576 4347
rect 4628 4312 4634 4364
rect 4970 4356 4978 4412
rect 5084 4370 5092 4422
rect 5034 4356 5092 4370
rect 4970 4347 5092 4356
rect 4974 4340 5092 4347
rect 4570 4301 4634 4312
rect 4566 4030 4630 4041
rect 4566 4013 4572 4030
rect 4466 4004 4572 4013
rect 4466 3948 4474 4004
rect 4530 3978 4572 4004
rect 4624 3978 4630 4030
rect 4530 3967 4630 3978
rect 4958 4004 5152 4022
rect 4530 3948 4598 3967
rect 4466 3939 4598 3948
rect 4958 3948 4978 4004
rect 5034 3970 5152 4004
rect 5034 3948 5036 3970
rect 4958 3918 5036 3948
rect 5088 3918 5152 3970
rect 4958 3902 5152 3918
rect 4958 3846 4978 3902
rect 5034 3852 5152 3902
rect 5034 3846 5036 3852
rect 4466 3805 4598 3809
rect 4466 3800 4630 3805
rect 4466 3744 4474 3800
rect 4530 3794 4630 3800
rect 4530 3744 4572 3794
rect 4466 3742 4572 3744
rect 4624 3742 4630 3794
rect 4466 3735 4630 3742
rect 4566 3731 4630 3735
rect 4958 3800 5036 3846
rect 5088 3800 5152 3852
rect 4958 3734 5152 3800
rect 4958 3698 5036 3734
rect 4958 3642 4978 3698
rect 5034 3682 5036 3698
rect 5088 3682 5152 3734
rect 5034 3642 5152 3682
rect 4958 3616 5152 3642
rect 4466 3596 4598 3605
rect 4466 3540 4474 3596
rect 4530 3569 4598 3596
rect 4958 3596 5036 3616
rect 4530 3558 4630 3569
rect 4530 3540 4572 3558
rect 4466 3531 4572 3540
rect 4566 3506 4572 3531
rect 4624 3506 4630 3558
rect 4958 3540 4978 3596
rect 5034 3564 5036 3596
rect 5088 3564 5152 3616
rect 5034 3540 5152 3564
rect 4958 3522 5152 3540
rect 4566 3495 4630 3506
<< via2 >>
rect 4726 11190 4782 11246
rect 5230 11224 5286 11246
rect 5230 11190 5270 11224
rect 5270 11190 5286 11224
rect 5230 11106 5286 11144
rect 5230 11088 5270 11106
rect 5270 11088 5286 11106
rect 4726 10986 4782 11042
rect 5230 10936 5270 10940
rect 5270 10936 5286 10940
rect 5230 10884 5286 10936
rect 3970 10782 4026 10838
rect 4726 10782 4782 10838
rect 4978 10782 5034 10838
rect 5230 10818 5270 10838
rect 5270 10818 5286 10838
rect 5230 10782 5286 10818
rect 4726 10374 4782 10430
rect 4978 10374 5034 10430
rect 5230 10418 5286 10430
rect 5230 10374 5270 10418
rect 5270 10374 5286 10418
rect 5230 10300 5286 10328
rect 5230 10272 5270 10300
rect 5270 10272 5286 10300
rect 4726 10170 4782 10226
rect 5230 10182 5286 10226
rect 5230 10170 5270 10182
rect 5270 10170 5286 10182
rect 4474 9966 4530 10022
rect 4726 9966 4782 10022
rect 4978 9966 5034 10022
rect 5230 10012 5270 10022
rect 5270 10012 5286 10022
rect 5230 9966 5286 10012
rect 4726 9660 4782 9716
rect 4978 9660 5034 9716
rect 5230 9612 5286 9614
rect 5230 9560 5270 9612
rect 5270 9560 5286 9612
rect 5230 9558 5286 9560
rect 5230 9494 5286 9512
rect 5230 9456 5270 9494
rect 5270 9456 5286 9494
rect 4726 9354 4782 9410
rect 5230 9376 5286 9410
rect 5230 9354 5270 9376
rect 5270 9354 5286 9376
rect 5230 9258 5286 9308
rect 5230 9252 5270 9258
rect 5270 9252 5286 9258
rect 4726 9150 4782 9206
rect 4978 9150 5034 9206
rect 4474 8844 4530 8900
rect 4726 8844 4782 8900
rect 4978 8742 5034 8798
rect 4978 8640 5034 8696
rect 4726 8538 4782 8594
rect 4978 8538 5034 8594
rect 4978 8436 5034 8492
rect 4222 8334 4278 8390
rect 4726 8334 4782 8390
rect 4726 8130 4782 8186
rect 4978 8130 5034 8186
rect 4474 8028 4530 8084
rect 4726 8028 4782 8084
rect 4978 7926 5034 7982
rect 5230 7926 5286 7982
rect 4474 7722 4530 7778
rect 4978 7824 5034 7880
rect 4978 7722 5034 7778
rect 4726 7620 4782 7676
rect 4978 7620 5034 7676
rect 4474 7518 4530 7574
rect 4474 7212 4530 7268
rect 4726 7212 4782 7268
rect 4978 7110 5034 7166
rect 4474 7008 4530 7064
rect 4978 7008 5034 7064
rect 4978 6906 5034 6962
rect 4978 6804 5034 6860
rect 4474 6702 4530 6758
rect 4222 6498 4278 6554
rect 4726 6498 4782 6554
rect 3970 6396 4026 6452
rect 4726 6294 4782 6350
rect 5230 6294 5286 6350
rect 3970 6192 4026 6248
rect 4222 6192 4278 6248
rect 5230 6192 5286 6248
rect 5230 6090 5286 6146
rect 4222 5886 4278 5942
rect 5230 5988 5286 6044
rect 4726 5886 4782 5942
rect 4726 5784 4782 5840
rect 5230 5784 5286 5840
rect 4474 5580 4530 5636
rect 4978 5530 5032 5534
rect 5032 5530 5034 5534
rect 4978 5478 5034 5530
rect 4474 5376 4530 5432
rect 4978 5412 5032 5432
rect 5032 5412 5034 5432
rect 4978 5376 5034 5412
rect 4978 5294 5032 5330
rect 5032 5294 5034 5330
rect 4978 5274 5034 5294
rect 4474 5070 4530 5126
rect 4726 5172 4782 5228
rect 4978 5176 5032 5228
rect 5032 5176 5034 5228
rect 4978 5172 5034 5176
rect 4474 4764 4530 4820
rect 4726 4764 4782 4820
rect 4978 4776 5034 4820
rect 4978 4764 5032 4776
rect 5032 4764 5034 4776
rect 5230 4764 5286 4820
rect 4474 4560 4530 4616
rect 4978 4606 5032 4616
rect 5032 4606 5034 4616
rect 4978 4560 5034 4606
rect 4978 4488 5032 4514
rect 5032 4488 5034 4514
rect 4978 4458 5034 4488
rect 4474 4356 4530 4412
rect 4978 4370 5032 4412
rect 5032 4370 5034 4412
rect 4978 4356 5034 4370
rect 4474 3948 4530 4004
rect 4978 3948 5034 4004
rect 4978 3846 5034 3902
rect 4474 3744 4530 3800
rect 4978 3642 5034 3698
rect 4474 3540 4530 3596
rect 4978 3540 5034 3596
<< metal3 >>
rect 4674 11246 4834 11254
rect 4674 11190 4726 11246
rect 4782 11190 4834 11246
rect 4674 11042 4834 11190
rect 4674 10986 4726 11042
rect 4782 10986 4834 11042
rect 3918 10838 4078 10846
rect 3918 10782 3970 10838
rect 4026 10782 4078 10838
rect 3918 6452 4078 10782
rect 4674 10838 4834 10986
rect 5178 11246 5338 11254
rect 5178 11190 5230 11246
rect 5286 11190 5338 11246
rect 5178 11144 5338 11190
rect 5178 11088 5230 11144
rect 5286 11088 5338 11144
rect 5178 10940 5338 11088
rect 5178 10884 5230 10940
rect 5286 10884 5338 10940
rect 4674 10782 4726 10838
rect 4782 10782 4834 10838
rect 4674 10774 4834 10782
rect 4926 10838 5086 10846
rect 4926 10782 4978 10838
rect 5034 10782 5086 10838
rect 4674 10430 4834 10438
rect 4674 10374 4726 10430
rect 4782 10374 4834 10430
rect 4674 10226 4834 10374
rect 4926 10430 5086 10782
rect 5178 10838 5338 10884
rect 5178 10782 5230 10838
rect 5286 10782 5338 10838
rect 5178 10774 5338 10782
rect 4926 10374 4978 10430
rect 5034 10374 5086 10430
rect 4926 10366 5086 10374
rect 5178 10430 5338 10438
rect 5178 10374 5230 10430
rect 5286 10374 5338 10430
rect 4674 10170 4726 10226
rect 4782 10170 4834 10226
rect 4422 10022 4582 10030
rect 4422 9966 4474 10022
rect 4530 9966 4582 10022
rect 4422 8900 4582 9966
rect 4674 10022 4834 10170
rect 5178 10328 5338 10374
rect 5178 10272 5230 10328
rect 5286 10272 5338 10328
rect 5178 10226 5338 10272
rect 5178 10170 5230 10226
rect 5286 10170 5338 10226
rect 4674 9966 4726 10022
rect 4782 9966 4834 10022
rect 4674 9958 4834 9966
rect 4926 10022 5086 10030
rect 4926 9966 4978 10022
rect 5034 9966 5086 10022
rect 4674 9716 4834 9724
rect 4674 9660 4726 9716
rect 4782 9660 4834 9716
rect 4674 9410 4834 9660
rect 4926 9716 5086 9966
rect 5178 10022 5338 10170
rect 5178 9966 5230 10022
rect 5286 9966 5338 10022
rect 5178 9958 5338 9966
rect 4926 9660 4978 9716
rect 5034 9660 5086 9716
rect 4926 9652 5086 9660
rect 4674 9354 4726 9410
rect 4782 9354 4834 9410
rect 4674 9206 4834 9354
rect 5178 9614 5338 9622
rect 5178 9558 5230 9614
rect 5286 9558 5338 9614
rect 5178 9512 5338 9558
rect 5178 9456 5230 9512
rect 5286 9456 5338 9512
rect 5178 9410 5338 9456
rect 5178 9354 5230 9410
rect 5286 9354 5338 9410
rect 5178 9308 5338 9354
rect 5178 9252 5230 9308
rect 5286 9252 5338 9308
rect 4674 9150 4726 9206
rect 4782 9150 4834 9206
rect 4674 9142 4834 9150
rect 4926 9206 5086 9214
rect 4926 9150 4978 9206
rect 5034 9150 5086 9206
rect 4422 8844 4474 8900
rect 4530 8844 4582 8900
rect 4422 8836 4582 8844
rect 4674 8900 4834 8908
rect 4674 8844 4726 8900
rect 4782 8844 4834 8900
rect 4674 8594 4834 8844
rect 4674 8538 4726 8594
rect 4782 8538 4834 8594
rect 4170 8390 4330 8398
rect 4170 8334 4222 8390
rect 4278 8334 4330 8390
rect 4170 6554 4330 8334
rect 4674 8390 4834 8538
rect 4674 8334 4726 8390
rect 4782 8334 4834 8390
rect 4674 8326 4834 8334
rect 4926 8798 5086 9150
rect 4926 8742 4978 8798
rect 5034 8742 5086 8798
rect 4926 8696 5086 8742
rect 4926 8640 4978 8696
rect 5034 8640 5086 8696
rect 4926 8594 5086 8640
rect 4926 8538 4978 8594
rect 5034 8538 5086 8594
rect 4926 8492 5086 8538
rect 4926 8436 4978 8492
rect 5034 8436 5086 8492
rect 4674 8186 4834 8194
rect 4674 8130 4726 8186
rect 4782 8130 4834 8186
rect 4422 8084 4582 8092
rect 4422 8028 4474 8084
rect 4530 8028 4582 8084
rect 4422 7778 4582 8028
rect 4674 8084 4834 8130
rect 4926 8186 5086 8436
rect 4926 8130 4978 8186
rect 5034 8130 5086 8186
rect 4926 8122 5086 8130
rect 4674 8028 4726 8084
rect 4782 8028 4834 8084
rect 4674 8020 4834 8028
rect 4422 7722 4474 7778
rect 4530 7722 4582 7778
rect 4422 7574 4582 7722
rect 4926 7982 5086 7990
rect 4926 7926 4978 7982
rect 5034 7926 5086 7982
rect 4926 7880 5086 7926
rect 5178 7982 5338 9252
rect 5178 7926 5230 7982
rect 5286 7926 5338 7982
rect 5178 7918 5338 7926
rect 4926 7824 4978 7880
rect 5034 7824 5086 7880
rect 4926 7778 5086 7824
rect 4926 7722 4978 7778
rect 5034 7722 5086 7778
rect 4422 7518 4474 7574
rect 4530 7518 4582 7574
rect 4422 7510 4582 7518
rect 4674 7676 4834 7684
rect 4674 7620 4726 7676
rect 4782 7620 4834 7676
rect 4170 6498 4222 6554
rect 4278 6498 4330 6554
rect 4170 6490 4330 6498
rect 4422 7268 4582 7276
rect 4422 7212 4474 7268
rect 4530 7212 4582 7268
rect 4422 7064 4582 7212
rect 4674 7268 4834 7620
rect 4926 7676 5086 7722
rect 4926 7620 4978 7676
rect 5034 7620 5086 7676
rect 4926 7612 5086 7620
rect 4674 7212 4726 7268
rect 4782 7212 4834 7268
rect 4674 7204 4834 7212
rect 4422 7008 4474 7064
rect 4530 7008 4582 7064
rect 4422 6758 4582 7008
rect 4422 6702 4474 6758
rect 4530 6702 4582 6758
rect 3918 6396 3970 6452
rect 4026 6396 4078 6452
rect 3918 6248 4078 6396
rect 3918 6192 3970 6248
rect 4026 6192 4078 6248
rect 3918 6184 4078 6192
rect 4170 6248 4330 6256
rect 4170 6192 4222 6248
rect 4278 6192 4330 6248
rect 4170 5942 4330 6192
rect 4170 5886 4222 5942
rect 4278 5886 4330 5942
rect 4170 5878 4330 5886
rect 4422 5636 4582 6702
rect 4926 7166 5086 7174
rect 4926 7110 4978 7166
rect 5034 7110 5086 7166
rect 4926 7064 5086 7110
rect 4926 7008 4978 7064
rect 5034 7008 5086 7064
rect 4926 6962 5086 7008
rect 4926 6906 4978 6962
rect 5034 6906 5086 6962
rect 4926 6860 5086 6906
rect 4926 6804 4978 6860
rect 5034 6804 5086 6860
rect 4674 6554 4834 6562
rect 4674 6498 4726 6554
rect 4782 6498 4834 6554
rect 4674 6350 4834 6498
rect 4674 6294 4726 6350
rect 4782 6294 4834 6350
rect 4674 6286 4834 6294
rect 4674 5942 4834 5950
rect 4674 5886 4726 5942
rect 4782 5886 4834 5942
rect 4674 5840 4834 5886
rect 4674 5784 4726 5840
rect 4782 5784 4834 5840
rect 4674 5776 4834 5784
rect 4422 5580 4474 5636
rect 4530 5580 4582 5636
rect 4422 5432 4582 5580
rect 4422 5376 4474 5432
rect 4530 5376 4582 5432
rect 4422 5126 4582 5376
rect 4926 5534 5086 6804
rect 5178 6350 5338 6358
rect 5178 6294 5230 6350
rect 5286 6294 5338 6350
rect 5178 6248 5338 6294
rect 5178 6192 5230 6248
rect 5286 6192 5338 6248
rect 5178 6146 5338 6192
rect 5178 6090 5230 6146
rect 5286 6090 5338 6146
rect 5178 6044 5338 6090
rect 5178 5988 5230 6044
rect 5286 5988 5338 6044
rect 5178 5980 5338 5988
rect 4926 5478 4978 5534
rect 5034 5478 5086 5534
rect 4926 5432 5086 5478
rect 4926 5376 4978 5432
rect 5034 5376 5086 5432
rect 4926 5330 5086 5376
rect 4926 5274 4978 5330
rect 5034 5274 5086 5330
rect 4422 5070 4474 5126
rect 4530 5070 4582 5126
rect 4422 5062 4582 5070
rect 4674 5228 4834 5236
rect 4674 5172 4726 5228
rect 4782 5172 4834 5228
rect 4422 4820 4582 4828
rect 4422 4764 4474 4820
rect 4530 4764 4582 4820
rect 4422 4616 4582 4764
rect 4674 4820 4834 5172
rect 4926 5228 5086 5274
rect 4926 5172 4978 5228
rect 5034 5172 5086 5228
rect 4926 5164 5086 5172
rect 5178 5840 5338 5848
rect 5178 5784 5230 5840
rect 5286 5784 5338 5840
rect 4674 4764 4726 4820
rect 4782 4764 4834 4820
rect 4674 4756 4834 4764
rect 4926 4820 5086 4828
rect 4926 4764 4978 4820
rect 5034 4764 5086 4820
rect 4422 4560 4474 4616
rect 4530 4560 4582 4616
rect 4422 4412 4582 4560
rect 4422 4356 4474 4412
rect 4530 4356 4582 4412
rect 4422 4004 4582 4356
rect 4422 3948 4474 4004
rect 4530 3948 4582 4004
rect 4422 3800 4582 3948
rect 4422 3744 4474 3800
rect 4530 3744 4582 3800
rect 4422 3596 4582 3744
rect 4422 3540 4474 3596
rect 4530 3540 4582 3596
rect 4422 3532 4582 3540
rect 4926 4616 5086 4764
rect 5178 4820 5338 5784
rect 5178 4764 5230 4820
rect 5286 4764 5338 4820
rect 5178 4756 5338 4764
rect 4926 4560 4978 4616
rect 5034 4560 5086 4616
rect 4926 4514 5086 4560
rect 4926 4458 4978 4514
rect 5034 4458 5086 4514
rect 4926 4412 5086 4458
rect 4926 4356 4978 4412
rect 5034 4356 5086 4412
rect 4926 4004 5086 4356
rect 4926 3948 4978 4004
rect 5034 3948 5086 4004
rect 4926 3902 5086 3948
rect 4926 3846 4978 3902
rect 5034 3846 5086 3902
rect 4926 3698 5086 3846
rect 4926 3642 4978 3698
rect 5034 3642 5086 3698
rect 4926 3596 5086 3642
rect 4926 3540 4978 3596
rect 5034 3540 5086 3596
rect 4926 3532 5086 3540
use XM1  XM1_0 ../Devices
timestamp 1691653953
transform 0 1 4634 -1 0 5380
box -403 -579 403 579
use XM2  XM2_0 ../Devices
timestamp 1691653953
transform 0 1 4634 -1 0 6992
box -403 -584 403 584
use XM3  XM3_0 ../Devices
timestamp 1691653953
transform 0 1 4872 -1 0 9410
box -403 -579 403 579
use XM4  XM4_0 ../Devices
timestamp 1691653953
transform 0 1 4634 -1 0 7798
box -403 -584 403 584
use XM5  XM5_0 ../Devices
timestamp 1691653953
transform 0 1 4872 -1 0 10216
box -403 -579 403 579
use XM6  XM6_0 ../Devices
timestamp 1691653953
transform 0 1 4872 -1 0 8604
box -403 -584 403 584
use XM7  XM7_0 ../Devices
timestamp 1691653954
transform 0 1 4872 -1 0 11022
box -403 -579 403 579
use XM8  XM8_0 ../Devices
timestamp 1691653954
transform 0 1 4634 -1 0 6186
box -403 -584 403 584
use XM9  XM9_0 ../Devices
timestamp 1691653954
transform 0 1 4634 -1 0 4574
box -403 -579 403 579
use XM10  XM10_0 ../Devices
timestamp 1691653954
transform 0 1 4634 -1 0 3768
box -403 -584 403 584
<< labels >>
rlabel via2 5006 7750 5006 7750 1 v1
rlabel via2 5006 7138 5006 7138 1 v0
rlabel via2 5006 8566 5006 8566 1 v2
rlabel metal2 4922 10402 4922 10402 1 v3
rlabel metal3 3998 6934 3998 6934 1 v4
<< end >>
