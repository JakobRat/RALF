** sch_path: /home/jakob/Documents/AutomatedLayoutGeneration/Circuits/Comparator/adc_comp_latch.sch
**.subckt adc_comp_latch VDD VSS clk inp inn comp_trig latch_qn latch_q
*.iopin VDD
*.iopin VSS
*.ipin clk
*.ipin inp
*.ipin inn
*.opin comp_trig
*.opin latch_qn
*.opin latch_q
x4 VDD VSS clk net1 adc_inverter
x5 VDD VSS net1 net2 adc_inverter
x3 comp_outp comp_outn VDD comp_trig VSS adc_nor
x2 comp_outp latch_qn VDD latch_q VSS comp_outn adc_nor_latch
x1 net2 net1 VDD comp_outp comp_outn inn inp VSS adc_comp
**.ends

* expanding   symbol:  adc_inverter.sym # of pins=4
** sym_path: /home/jakob/Documents/AutomatedLayoutGeneration/Circuits/Comparator/adc_inverter.sym
** sch_path: /home/jakob/Documents/AutomatedLayoutGeneration/Circuits/Comparator/adc_inverter.sch
.subckt adc_inverter VDD VSS in out
*.iopin VDD
*.iopin VSS
*.ipin in
*.opin out
XM2 out in VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=0.84 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM1 out in VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  adc_nor.sym # of pins=5
** sym_path: /home/jakob/Documents/AutomatedLayoutGeneration/Circuits/Comparator/adc_nor.sym
** sch_path: /home/jakob/Documents/AutomatedLayoutGeneration/Circuits/Comparator/adc_nor.sch
.subckt adc_nor b a VDD q VSS
*.iopin VDD
*.iopin VSS
*.ipin b
*.ipin a
*.opin q
XM5 q b VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM6 q a VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM1 q b net1 VDD sky130_fd_pr__pfet_01v8 L=0.15 W=0.8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM2 q a net2 VDD sky130_fd_pr__pfet_01v8 L=0.15 W=0.8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM3 net2 b VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=0.8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM4 net1 a VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=0.8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  adc_nor_latch.sym # of pins=6
** sym_path: /home/jakob/Documents/AutomatedLayoutGeneration/Circuits/Comparator/adc_nor_latch.sym
** sch_path: /home/jakob/Documents/AutomatedLayoutGeneration/Circuits/Comparator/adc_nor_latch.sch
.subckt adc_nor_latch s qn VDD q VSS r
*.iopin VDD
*.iopin VSS
*.ipin s
*.ipin r
*.opin q
*.opin qn
x1 q s VDD qn VSS adc_nor
x2 qn r VDD q VSS adc_nor
.ends


* expanding   symbol:
*+  /home/jakob/Documents/AutomatedLayoutGeneration/Circuits/Comparator/adc_comp.sym # of pins=8
** sym_path: /home/jakob/Documents/AutomatedLayoutGeneration/Circuits/Comparator/adc_comp.sym
** sch_path: /home/jakob/Documents/AutomatedLayoutGeneration/Circuits/Comparator/adc_comp.sch
.subckt adc_comp clk nclk VPWR outp outn inn inp VGND
*.iopin VPWR
*.iopin VGND
*.ipin clk
*.ipin nclk
*.ipin inp
*.ipin inn
*.opin outp
*.opin outn
XC1 on VGND sky130_fd_pr__cap_mim_m3_1 W=18.9 L=5.1 MF=1 m=1
XC2 op VGND sky130_fd_pr__cap_mim_m3_1 W=18.9 L=5.1 MF=1 m=1
x1 clk nclk VPWR on op inn inp VGND DiffAmp
x2 clk nclk VPWR outp_nb op on outn_nb VGND Comp
x3 VPWR VGND outp_nb outp adc_comp_buffer
x4 VPWR VGND outn_nb outn adc_comp_buffer
.ends


* expanding   symbol:
*+  /home/jakob/Documents/AutomatedLayoutGeneration/Circuits/Comparator/DiffAmp.sym # of pins=8
** sym_path: /home/jakob/Documents/AutomatedLayoutGeneration/Circuits/Comparator/DiffAmp.sym
** sch_path: /home/jakob/Documents/AutomatedLayoutGeneration/Circuits/Comparator/DiffAmp.sch
.subckt DiffAmp clk nclk VPWR outn outp inn inp VGND
*.iopin VPWR
*.iopin VGND
*.ipin clk
*.ipin nclk
*.ipin inp
*.ipin inn
*.opin outn
*.opin outp
XM3 outn inp in_stage_net1 VGND sky130_fd_pr__nfet_01v8 L=0.15 W=8 nf=4 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM4 outp inn in_stage_net1 VGND sky130_fd_pr__nfet_01v8 L=0.15 W=8 nf=4 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM5 in_stage_net1 clk VGND VGND sky130_fd_pr__nfet_01v8 L=0.15 W=4 nf=8 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM2 outp clk VPWR VPWR sky130_fd_pr__pfet_01v8 L=0.15 W=2 nf=4 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM1 outn clk VPWR VPWR sky130_fd_pr__pfet_01v8 L=0.15 W=2 nf=4 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  /home/jakob/Documents/AutomatedLayoutGeneration/Circuits/Comparator/Comp.sym
*+ # of pins=8
** sym_path: /home/jakob/Documents/AutomatedLayoutGeneration/Circuits/Comparator/Comp.sym
** sch_path: /home/jakob/Documents/AutomatedLayoutGeneration/Circuits/Comparator/Comp.sch
.subckt Comp clk nclk VPWR outp inp inn outn VGND
*.opin outp
*.opin outn
*.iopin VPWR
*.ipin clk
*.ipin nclk
*.iopin VGND
*.ipin inp
*.ipin inn
XM6 in_stage_net2 outp VPWR VPWR sky130_fd_pr__pfet_01v8 L=0.15 W=4 nf=2 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM7 in_stage_net3 outn VPWR VPWR sky130_fd_pr__pfet_01v8 L=0.15 W=4 nf=2 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM8 outn inn in_stage_net2 VPWR sky130_fd_pr__pfet_01v8 L=0.15 W=4 nf=2 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM9 outp inp in_stage_net3 VPWR sky130_fd_pr__pfet_01v8 L=0.15 W=4 nf=2 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM10 outn outp VGND VGND sky130_fd_pr__nfet_01v8 L=0.15 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM11 outn nclk VGND VGND sky130_fd_pr__nfet_01v8 L=0.15 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM12 outp nclk VGND VGND sky130_fd_pr__nfet_01v8 L=0.15 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM13 outp outn VGND VGND sky130_fd_pr__nfet_01v8 L=0.15 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  adc_comp_buffer.sym # of pins=4
** sym_path: /home/jakob/Documents/AutomatedLayoutGeneration/Circuits/Comparator/adc_comp_buffer.sym
** sch_path: /home/jakob/Documents/AutomatedLayoutGeneration/Circuits/Comparator/adc_comp_buffer.sch
.subckt adc_comp_buffer VDD VSS in out
*.iopin VDD
*.iopin VSS
*.ipin in
*.opin out
XM5 buf_mid in VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM1 buf_mid in VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM2 out buf_mid VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=2 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM6 out buf_mid VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
.ends

.end
