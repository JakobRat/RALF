magic
tech sky130A
timestamp 1702577692
<< checkpaint >>
rect -1187 -1104 1187 1104
<< pwell >>
rect -557 -474 557 474
<< psubdiff >>
rect -539 439 539 456
rect -539 -439 -522 439
rect 522 -439 539 439
rect -539 -456 -491 -439
rect 491 -456 539 -439
<< psubdiffcont >>
rect -491 -456 491 -439
<< xpolycontact >>
rect -474 175 -439 391
rect -474 -391 -439 -175
rect -391 175 -356 391
rect -391 -391 -356 -175
rect -308 175 -273 391
rect -308 -391 -273 -175
rect -225 175 -190 391
rect -225 -391 -190 -175
rect -142 175 -107 391
rect -142 -391 -107 -175
rect -59 175 -24 391
rect -59 -391 -24 -175
rect 24 175 59 391
rect 24 -391 59 -175
rect 107 175 142 391
rect 107 -391 142 -175
rect 190 175 225 391
rect 190 -391 225 -175
rect 273 175 308 391
rect 273 -391 308 -175
rect 356 175 391 391
rect 356 -391 391 -175
rect 439 175 474 391
rect 439 -391 474 -175
<< xpolyres >>
rect -474 -175 -439 175
rect -391 -175 -356 175
rect -308 -175 -273 175
rect -225 -175 -190 175
rect -142 -175 -107 175
rect -59 -175 -24 175
rect 24 -175 59 175
rect 107 -175 142 175
rect 190 -175 225 175
rect 273 -175 308 175
rect 356 -175 391 175
rect 439 -175 474 175
<< locali >>
rect -499 -456 -491 -439
rect 491 -456 499 -439
<< res0p35 >>
rect -475 -176 -438 176
rect -392 -176 -355 176
rect -309 -176 -272 176
rect -226 -176 -189 176
rect -143 -176 -106 176
rect -60 -176 -23 176
rect 23 -176 60 176
rect 106 -176 143 176
rect 189 -176 226 176
rect 272 -176 309 176
rect 355 -176 392 176
rect 438 -176 475 176
<< properties >>
string FIXED_BBOX -530 -447 530 447
<< end >>
