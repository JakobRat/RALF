magic
tech sky130A
magscale 1 2
timestamp 1702541238
<< checkpaint >>
rect -1556 -2244 1556 2244
<< nwell >>
rect -296 -984 296 984
<< pmos >>
rect -100 -836 100 764
<< pdiff >>
rect -158 752 -100 764
rect -158 -824 -146 752
rect -112 -824 -100 752
rect -158 -836 -100 -824
rect 100 752 158 764
rect 100 -824 112 752
rect 146 -824 158 752
rect 100 -836 158 -824
<< pdiffc >>
rect -146 -824 -112 752
rect 112 -824 146 752
<< nsubdiff >>
rect -260 914 260 948
rect -260 -914 -226 914
rect 226 -914 260 914
rect -260 -948 -164 -914
rect 164 -948 260 -914
<< nsubdiffcont >>
rect -164 -948 164 -914
<< poly >>
rect -100 845 100 861
rect -100 811 -84 845
rect 84 811 100 845
rect -100 764 100 811
rect -100 -862 100 -836
<< polycont >>
rect -84 811 84 845
<< locali >>
rect -260 914 260 948
rect -260 -914 -226 914
rect -100 811 -84 845
rect 84 811 100 845
rect -146 752 -112 768
rect -146 -840 -112 -824
rect 112 752 146 768
rect 112 -840 146 -824
rect 226 -914 260 914
rect -260 -948 -164 -914
rect 164 -948 260 -914
<< properties >>
string FIXED_BBOX -243 -931 243 931
<< end >>
