magic
tech sky130A
magscale 1 2
timestamp 1701085297
<< checkpaint >>
rect -1261 2109 2109 2333
rect -1261 2052 2667 2109
rect -1261 1797 3225 2052
rect -1685 -1260 3225 1797
rect -1685 -1261 2667 -1260
rect -1685 -1797 1685 -1261
use XDL_XM3_XM4  XDL_XM3_XM4_0 ~/Documents/RALF/Magic/Devices
timestamp 1701085217
transform 1 0 424 0 1 536
box -425 -537 425 537
use XDP_XM1_XM2  XDP_XM1_XM2_0 ~/Documents/RALF/Magic/Devices
timestamp 1701085217
transform 0 -1 1128 1 0 424
box -425 -279 425 279
use XM5  XM5_0 ~/Documents/RALF/Magic/Devices
timestamp 1701085217
transform 0 1 1686 -1 0 396
box -396 -279 396 279
<< end >>
