** sch_path: /home/jakob/Documents/AutomatedLayoutGeneration/Circuits/CrossCoupledPair/CCP.sch
**.subckt CCP Vd1 Vd2 Vs2 Vs1 Vb
*.iopin Vd1
*.iopin Vd2
*.iopin Vs2
*.iopin Vs1
*.iopin Vb
XM1 Vd1 Vd2 Vs Vb sky130_fd_pr__nfet_01v8 L=0.5 W=20 nf=10 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM2 Vd2 Vd1 Vs Vb sky130_fd_pr__nfet_01v8 L=0.5 W=20 nf=10 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
**.ends
.end