magic
tech sky130A
magscale 1 2
timestamp 1702630323
<< checkpaint >>
rect 1485 3314 4597 3415
rect 369 1997 4597 3314
rect -1556 1539 4597 1997
rect -1685 -579 4597 1539
rect -1685 -1539 1685 -579
rect -1556 -1997 1556 -1539
use XDL_XM3_XM4  XDL_XM3_XM4_0 ~/Documents/RALF/Magic/Devices
timestamp 1702630323
transform -1 0 3041 0 -1 1418
box -296 -737 296 737
use XDP_XM1_XM2  XDP_XM1_XM2_0 ~/Documents/RALF/Magic/Devices
timestamp 1702630323
transform 0 1 2466 -1 0 1434
box -425 -279 425 279
use XM5  XM5_0 ~/Documents/RALF/Magic/Devices
timestamp 1702630323
transform 0 -1 1908 1 0 1658
box -396 -279 396 279
<< end >>
