magic
tech sky130A
magscale 1 2
timestamp 1702977096
<< checkpaint >>
rect -1656 -2439 1656 2439
<< pwell >>
rect -396 -1179 396 1179
<< nmos >>
rect -200 -1031 200 969
<< ndiff >>
rect -258 957 -200 969
rect -258 -1019 -246 957
rect -212 -1019 -200 957
rect -258 -1031 -200 -1019
rect 200 957 258 969
rect 200 -1019 212 957
rect 246 -1019 258 957
rect 200 -1031 258 -1019
<< ndiffc >>
rect -246 -1019 -212 957
rect 212 -1019 246 957
<< psubdiff >>
rect -360 1109 360 1143
rect -360 -1109 -326 1109
rect 326 -1109 360 1109
rect -360 -1143 -264 -1109
rect 264 -1143 360 -1109
<< psubdiffcont >>
rect -264 -1143 264 -1109
<< poly >>
rect -200 1041 200 1057
rect -200 1007 -184 1041
rect 184 1007 200 1041
rect -200 969 200 1007
rect -200 -1057 200 -1031
<< polycont >>
rect -184 1007 184 1041
<< locali >>
rect -360 1109 360 1143
rect -360 -1109 -326 1109
rect -200 1007 -184 1041
rect 184 1007 200 1041
rect -246 957 -212 973
rect -246 -1035 -212 -1019
rect 212 957 246 973
rect 212 -1035 246 -1019
rect 326 -1109 360 1109
rect -360 -1143 -264 -1109
rect 264 -1143 360 -1109
<< properties >>
string FIXED_BBOX -343 -1126 343 1126
<< end >>
