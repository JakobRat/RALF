magic
tech sky130A
magscale 1 2
timestamp 1701937757
<< checkpaint >>
rect -526 4613 3068 4617
rect -526 4025 4300 4613
rect -1260 3067 4300 4025
rect -1261 2109 4509 3067
rect -1261 2033 4617 2109
rect -1876 -1261 4617 2033
rect -1876 -2033 1876 -1261
use XCCP_XM3_XM4_x1  XCCP_XM3_XM4_x1_0 ~/Documents/RALF/Magic/Devices
timestamp 1701937427
transform -1 0 2103 0 -1 1270
box -296 -537 296 537
use XCCP_XM3_XM4_x2  XCCP_XM3_XM4_x2_0 ~/Documents/RALF/Magic/Devices
timestamp 1701937427
transform -1 0 295 0 -1 1270
box -296 -537 296 537
use XCCP_XM3_XM4_x3  XCCP_XM3_XM4_x3_0 ~/Documents/RALF/Magic/Devices
timestamp 1701937428
transform 0 -1 1271 1 0 3061
box -296 -537 296 537
use XDP_XM1_XM2_x1  XDP_XM1_XM2_x1_0 ~/Documents/RALF/Magic/Devices
timestamp 1701937427
transform 1 0 2824 0 1 1328
box -425 -479 425 479
use XDP_XM1_XM2_x2  XDP_XM1_XM2_x2_0 ~/Documents/RALF/Magic/Devices
timestamp 1701937427
transform 1 0 1016 0 1 1328
box -425 -479 425 479
use XDP_XM1_XM2_x3  XDP_XM1_XM2_x3_0 ~/Documents/RALF/Magic/Devices
timestamp 1701937428
transform 0 1 1329 -1 0 2340
box -425 -479 425 479
use XM5_x1  XM5_x1_0 ~/Documents/RALF/Magic/Devices
timestamp 1701937427
transform 0 1 2878 -1 0 424
box -425 -479 425 479
use XM5_x2  XM5_x2_0 ~/Documents/RALF/Magic/Devices
timestamp 1701937427
transform 0 1 1070 -1 0 424
box -425 -479 425 479
use XM5_x3  XM5_x3_0 ~/Documents/RALF/Magic/Devices
timestamp 1701937428
transform -1 0 425 0 -1 2286
box -425 -479 425 479
use XRSTR_0  XRSTR_0_0 ~/Documents/RALF/Magic/Devices
timestamp 1701937426
transform 1 0 2424 0 1 2580
box -616 -773 616 773
<< end >>
