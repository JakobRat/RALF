magic
tech sky130A
magscale 1 2
timestamp 1701181053
<< checkpaint >>
rect -1685 -1797 1685 1797
<< nwell >>
rect -425 -537 425 537
<< pmos >>
rect -229 118 -29 318
rect 29 118 229 318
rect -229 -318 -29 -118
rect 29 -318 229 -118
<< pdiff >>
rect -287 306 -229 318
rect -287 130 -275 306
rect -241 130 -229 306
rect -287 118 -229 130
rect -29 306 29 318
rect -29 130 -17 306
rect 17 130 29 306
rect -29 118 29 130
rect 229 306 287 318
rect 229 130 241 306
rect 275 130 287 306
rect 229 118 287 130
rect -287 -130 -229 -118
rect -287 -306 -275 -130
rect -241 -306 -229 -130
rect -287 -318 -229 -306
rect -29 -130 29 -118
rect -29 -306 -17 -130
rect 17 -306 29 -130
rect -29 -318 29 -306
rect 229 -130 287 -118
rect 229 -306 241 -130
rect 275 -306 287 -130
rect 229 -318 287 -306
<< pdiffc >>
rect -275 130 -241 306
rect -17 130 17 306
rect 241 130 275 306
rect -275 -306 -241 -130
rect -17 -306 17 -130
rect 241 -306 275 -130
<< nsubdiff >>
rect -389 467 389 501
rect -389 -467 -355 467
rect 355 -467 389 467
rect -389 -501 -293 -467
rect 293 -501 389 -467
<< nsubdiffcont >>
rect -293 -501 293 -467
<< poly >>
rect -229 399 -29 415
rect -229 365 -213 399
rect -45 365 -29 399
rect -229 318 -29 365
rect 29 399 229 415
rect 29 365 45 399
rect 213 365 229 399
rect 29 318 229 365
rect -229 71 -29 118
rect -229 37 -213 71
rect -45 37 -29 71
rect -229 21 -29 37
rect 29 71 229 118
rect 29 37 45 71
rect 213 37 229 71
rect 29 21 229 37
rect -229 -37 -29 -21
rect -229 -71 -213 -37
rect -45 -71 -29 -37
rect -229 -118 -29 -71
rect 29 -37 229 -21
rect 29 -71 45 -37
rect 213 -71 229 -37
rect 29 -118 229 -71
rect -229 -365 -29 -318
rect -229 -399 -213 -365
rect -45 -399 -29 -365
rect -229 -415 -29 -399
rect 29 -365 229 -318
rect 29 -399 45 -365
rect 213 -399 229 -365
rect 29 -415 229 -399
<< polycont >>
rect -213 365 -45 399
rect 45 365 213 399
rect -213 37 -45 71
rect 45 37 213 71
rect -213 -71 -45 -37
rect 45 -71 213 -37
rect -213 -399 -45 -365
rect 45 -399 213 -365
<< locali >>
rect -389 467 389 501
rect -389 -467 -355 467
rect -229 365 -213 399
rect -45 365 -29 399
rect 29 365 45 399
rect 213 365 229 399
rect -275 306 -241 322
rect -275 114 -241 130
rect -17 306 17 322
rect -17 114 17 130
rect 241 306 275 322
rect 241 114 275 130
rect -229 37 -213 71
rect -45 37 -29 71
rect 29 37 45 71
rect 213 37 229 71
rect -229 -71 -213 -37
rect -45 -71 -29 -37
rect 29 -71 45 -37
rect 213 -71 229 -37
rect -275 -130 -241 -114
rect -275 -322 -241 -306
rect -17 -130 17 -114
rect -17 -322 17 -306
rect 241 -130 275 -114
rect 241 -322 275 -306
rect -229 -399 -213 -365
rect -45 -399 -29 -365
rect 29 -399 45 -365
rect 213 -399 229 -365
rect 355 -467 389 467
rect -389 -501 -293 -467
rect 293 -501 389 -467
<< properties >>
string FIXED_BBOX -372 -484 372 484
<< end >>
